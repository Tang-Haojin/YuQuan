module dual_AsyncQueueSink_5( 
  input         clock, 
  input         reset, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [19:0] io_deq_bits_a, 
  output [19:0] io_deq_bits_b, 
  output [19:0] io_deq_bits_c, 
  output [19:0] io_deq_bits_d, 
  output [19:0] io_deq_bits_e, 
  input  [19:0] io_async_mem_0_a, 
  input  [19:0] io_async_mem_0_b, 
  input  [19:0] io_async_mem_0_c, 
  input  [19:0] io_async_mem_0_d, 
  input  [19:0] io_async_mem_0_e, 
  output        io_async_ridx, 
  input         io_async_widx, 
  output        io_async_safe_ridx_valid, 
  input         io_async_safe_widx_valid, 
  input         io_async_safe_source_reset_n, 
  output        io_async_safe_sink_reset_n 
);
  wire  ridx_bin_clock; 
  wire  ridx_bin_reset; 
  wire  ridx_bin_io_d; 
  wire  ridx_bin_io_q; 
  wire  ridx_bin_io_en; 
  wire  widx_gray_clock; 
  wire  widx_gray_reset; 
  wire  widx_gray_io_d; 
  wire  widx_gray_io_q; 
  wire  deq_bits_reg_clock; 
  wire [99:0] deq_bits_reg_io_d; 
  wire [99:0] deq_bits_reg_io_q; 
  wire  valid_reg_clock; 
  wire  valid_reg_reset; 
  wire  valid_reg_io_d; 
  wire  valid_reg_io_q; 
  wire  valid_reg_io_en; 
  wire  ridx_gray_clock; 
  wire  ridx_gray_reset; 
  wire  ridx_gray_io_d; 
  wire  ridx_gray_io_q; 
  wire  ridx_gray_io_en; 
  wire  AsyncValidSync_clock; 
  wire  AsyncValidSync_reset; 
  wire  AsyncValidSync_io_in; 
  wire  AsyncValidSync_io_out; 
  wire  AsyncValidSync_1_clock; 
  wire  AsyncValidSync_1_reset; 
  wire  AsyncValidSync_1_io_in; 
  wire  AsyncValidSync_1_io_out; 
  wire  AsyncValidSync_2_clock; 
  wire  AsyncValidSync_2_reset; 
  wire  AsyncValidSync_2_io_in; 
  wire  AsyncValidSync_2_io_out; 
  wire  AsyncResetRegVec_w1_i0_clock; 
  wire  AsyncResetRegVec_w1_i0_reset; 
  wire  AsyncResetRegVec_w1_i0_io_d; 
  wire  AsyncResetRegVec_w1_i0_io_q; 
  wire  AsyncResetRegVec_w1_i0_io_en; 
  wire  _T; 
  wire  source_ready; 
  wire  _T_1; 
  wire  _T_4; 
  wire  ridx; 
  wire  widx; 
  wire  _T_7; 
  wire  valid; 
  wire [19:0] deq_bits_nxt_a; 
  wire [19:0] deq_bits_nxt_b; 
  wire [19:0] deq_bits_nxt_c; 
  wire [19:0] deq_bits_nxt_d; 
  wire [19:0] deq_bits_nxt_e; 
  wire [39:0] _T_8; 
  wire [59:0] _T_10; 
  wire [99:0] _T_13; 
  wire  valid_reg_1; 
  wire  _T_21; 
  dual_AsyncResetRegVec_w1_i0 ridx_bin ( 
    .clock(ridx_bin_clock),
    .reset(ridx_bin_reset),
    .io_d(ridx_bin_io_d),
    .io_q(ridx_bin_io_q),
    .io_en(ridx_bin_io_en)
  );
  dual_AsyncResetSynchronizerShiftReg_w1_d3_i0 widx_gray ( 
    .clock(widx_gray_clock),
    .reset(widx_gray_reset),
    .io_d(widx_gray_io_d),
    .io_q(widx_gray_io_q)
  );
  dual_SynchronizerShiftReg_w100_d1 deq_bits_reg ( 
    .clock(deq_bits_reg_clock),
    .io_d(deq_bits_reg_io_d),
    .io_q(deq_bits_reg_io_q)
  );
  dual_AsyncResetRegVec_w1_i0 valid_reg ( 
    .clock(valid_reg_clock),
    .reset(valid_reg_reset),
    .io_d(valid_reg_io_d),
    .io_q(valid_reg_io_q),
    .io_en(valid_reg_io_en)
  );
  dual_AsyncResetRegVec_w1_i0 ridx_gray ( 
    .clock(ridx_gray_clock),
    .reset(ridx_gray_reset),
    .io_d(ridx_gray_io_d),
    .io_q(ridx_gray_io_q),
    .io_en(ridx_gray_io_en)
  );
  dual_AsyncValidSync AsyncValidSync ( 
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_in(AsyncValidSync_io_in),
    .io_out(AsyncValidSync_io_out)
  );
  dual_AsyncValidSync_1 AsyncValidSync_1 ( 
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  dual_AsyncValidSync_2 AsyncValidSync_2 ( 
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  dual_AsyncResetRegVec_w1_i0 AsyncResetRegVec_w1_i0 ( 
    .clock(AsyncResetRegVec_w1_i0_clock),
    .reset(AsyncResetRegVec_w1_i0_reset),
    .io_d(AsyncResetRegVec_w1_i0_io_d),
    .io_q(AsyncResetRegVec_w1_i0_io_q),
    .io_en(AsyncResetRegVec_w1_i0_io_en)
  );
  assign _T = io_deq_ready & io_deq_valid; 
  assign source_ready = AsyncValidSync_2_io_out; 
  assign _T_1 = source_ready == 1'h0; 
  assign _T_4 = ridx_bin_io_q + _T; 
  assign ridx = _T_1 ? 1'h0 : _T_4; 
  assign widx = widx_gray_io_q; 
  assign _T_7 = ridx != widx; 
  assign valid = source_ready & _T_7; 
  assign deq_bits_nxt_a = valid ? io_async_mem_0_a : io_deq_bits_a; 
  assign deq_bits_nxt_b = valid ? io_async_mem_0_b : io_deq_bits_b; 
  assign deq_bits_nxt_c = valid ? io_async_mem_0_c : io_deq_bits_c; 
  assign deq_bits_nxt_d = valid ? io_async_mem_0_d : io_deq_bits_d; 
  assign deq_bits_nxt_e = valid ? io_async_mem_0_e : io_deq_bits_e; 
  assign _T_8 = {deq_bits_nxt_d,deq_bits_nxt_e}; 
  assign _T_10 = {deq_bits_nxt_a,deq_bits_nxt_b,deq_bits_nxt_c}; 
  assign _T_13 = deq_bits_reg_io_q; 
  assign valid_reg_1 = valid_reg_io_q; 
  assign _T_21 = io_async_safe_source_reset_n == 1'h0; 
  assign io_deq_valid = valid_reg_1 & source_ready; 
  assign io_deq_bits_a = _T_13[99:80]; 
  assign io_deq_bits_b = _T_13[79:60]; 
  assign io_deq_bits_c = _T_13[59:40]; 
  assign io_deq_bits_d = _T_13[39:20]; 
  assign io_deq_bits_e = _T_13[19:0]; 
  assign io_async_ridx = ridx_gray_io_q; 
  assign io_async_safe_ridx_valid = AsyncValidSync_io_out; 
  assign io_async_safe_sink_reset_n = reset == 1'h0; 
  assign ridx_bin_clock = clock; 
  assign ridx_bin_reset = reset; 
  assign ridx_bin_io_d = _T_1 ? 1'h0 : _T_4; 
  assign ridx_bin_io_en = 1'h1; 
  assign widx_gray_clock = clock; 
  assign widx_gray_reset = reset; 
  assign widx_gray_io_d = io_async_widx; 
  assign deq_bits_reg_clock = clock; 
  assign deq_bits_reg_io_d = {_T_10,_T_8}; 
  assign valid_reg_clock = clock; 
  assign valid_reg_reset = reset; 
  assign valid_reg_io_d = source_ready & _T_7; 
  assign valid_reg_io_en = 1'h1; 
  assign ridx_gray_clock = clock; 
  assign ridx_gray_reset = reset; 
  assign ridx_gray_io_d = _T_1 ? 1'h0 : _T_4; 
  assign ridx_gray_io_en = 1'h1; 
  assign AsyncValidSync_clock = clock; 
  assign AsyncValidSync_reset = reset | _T_21; 
  assign AsyncValidSync_io_in = 1'h1; 
  assign AsyncValidSync_1_clock = clock; 
  assign AsyncValidSync_1_reset = reset | _T_21; 
  assign AsyncValidSync_1_io_in = io_async_safe_widx_valid; 
  assign AsyncValidSync_2_clock = clock; 
  assign AsyncValidSync_2_reset = reset; 
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out; 
  assign AsyncResetRegVec_w1_i0_clock = clock; 
  assign AsyncResetRegVec_w1_i0_reset = reset; 
  assign AsyncResetRegVec_w1_i0_io_d = io_async_widx == io_async_ridx; 
  assign AsyncResetRegVec_w1_i0_io_en = 1'h1; 
endmodule
module dual_AsyncQueueSink( 
  input         clock, 
  input         reset, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [31:0] io_deq_bits, 
  input  [31:0] io_async_mem_0, 
  input  [31:0] io_async_mem_1, 
  input  [31:0] io_async_mem_2, 
  input  [31:0] io_async_mem_3, 
  input  [31:0] io_async_mem_4, 
  input  [31:0] io_async_mem_5, 
  input  [31:0] io_async_mem_6, 
  input  [31:0] io_async_mem_7, 
  output [3:0]  io_async_ridx, 
  input  [3:0]  io_async_widx, 
  output        io_async_safe_ridx_valid, 
  input         io_async_safe_widx_valid, 
  input         io_async_safe_source_reset_n, 
  output        io_async_safe_sink_reset_n 
);
  wire  ridx_bin_clock; 
  wire  ridx_bin_reset; 
  wire [3:0] ridx_bin_io_d; 
  wire [3:0] ridx_bin_io_q; 
  wire  ridx_bin_io_en; 
  wire  widx_gray_clock; 
  wire  widx_gray_reset; 
  wire [3:0] widx_gray_io_d; 
  wire [3:0] widx_gray_io_q; 
  wire  deq_bits_reg_clock; 
  wire [31:0] deq_bits_reg_io_d; 
  wire [31:0] deq_bits_reg_io_q; 
  wire  valid_reg_clock; 
  wire  valid_reg_reset; 
  wire  valid_reg_io_d; 
  wire  valid_reg_io_q; 
  wire  valid_reg_io_en; 
  wire  ridx_gray_clock; 
  wire  ridx_gray_reset; 
  wire [3:0] ridx_gray_io_d; 
  wire [3:0] ridx_gray_io_q; 
  wire  ridx_gray_io_en; 
  wire  AsyncValidSync_clock; 
  wire  AsyncValidSync_reset; 
  wire  AsyncValidSync_io_in; 
  wire  AsyncValidSync_io_out; 
  wire  AsyncValidSync_1_clock; 
  wire  AsyncValidSync_1_reset; 
  wire  AsyncValidSync_1_io_in; 
  wire  AsyncValidSync_1_io_out; 
  wire  AsyncValidSync_2_clock; 
  wire  AsyncValidSync_2_reset; 
  wire  AsyncValidSync_2_io_in; 
  wire  AsyncValidSync_2_io_out; 
  wire  AsyncResetRegVec_w1_i0_clock; 
  wire  AsyncResetRegVec_w1_i0_reset; 
  wire  AsyncResetRegVec_w1_i0_io_d; 
  wire  AsyncResetRegVec_w1_i0_io_q; 
  wire  AsyncResetRegVec_w1_i0_io_en; 
  wire  _T; 
  wire  source_ready; 
  wire  _T_1; 
  wire [3:0] _GEN_8; 
  wire [3:0] _T_4; 
  wire [3:0] _T_5; 
  wire [2:0] _T_6; 
  wire [3:0] _GEN_9; 
  wire [3:0] ridx; 
  wire [3:0] widx; 
  wire  _T_7; 
  wire  valid; 
  wire [2:0] _T_8; 
  wire  _T_9; 
  wire [2:0] _T_10; 
  wire [2:0] index; 
  wire [31:0] _GEN_1; 
  wire [31:0] _GEN_2; 
  wire [31:0] _GEN_3; 
  wire [31:0] _GEN_4; 
  wire [31:0] _GEN_5; 
  wire [31:0] _GEN_6; 
  wire [31:0] _GEN_7; 
  wire  valid_reg_1; 
  wire  _T_14; 
  dual_AsyncResetRegVec_w4_i0 ridx_bin ( 
    .clock(ridx_bin_clock),
    .reset(ridx_bin_reset),
    .io_d(ridx_bin_io_d),
    .io_q(ridx_bin_io_q),
    .io_en(ridx_bin_io_en)
  );
  dual_AsyncResetSynchronizerShiftReg_w4_d3_i0 widx_gray ( 
    .clock(widx_gray_clock),
    .reset(widx_gray_reset),
    .io_d(widx_gray_io_d),
    .io_q(widx_gray_io_q)
  );
  dual_SynchronizerShiftReg_w32_d1 deq_bits_reg ( 
    .clock(deq_bits_reg_clock),
    .io_d(deq_bits_reg_io_d),
    .io_q(deq_bits_reg_io_q)
  );
  dual_AsyncResetRegVec_w1_i0 valid_reg ( 
    .clock(valid_reg_clock),
    .reset(valid_reg_reset),
    .io_d(valid_reg_io_d),
    .io_q(valid_reg_io_q),
    .io_en(valid_reg_io_en)
  );
  dual_AsyncResetRegVec_w4_i0 ridx_gray ( 
    .clock(ridx_gray_clock),
    .reset(ridx_gray_reset),
    .io_d(ridx_gray_io_d),
    .io_q(ridx_gray_io_q),
    .io_en(ridx_gray_io_en)
  );
  dual_AsyncValidSync AsyncValidSync ( 
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_in(AsyncValidSync_io_in),
    .io_out(AsyncValidSync_io_out)
  );
  dual_AsyncValidSync_1 AsyncValidSync_1 ( 
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  dual_AsyncValidSync_2 AsyncValidSync_2 ( 
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  dual_AsyncResetRegVec_w1_i0 AsyncResetRegVec_w1_i0 ( 
    .clock(AsyncResetRegVec_w1_i0_clock),
    .reset(AsyncResetRegVec_w1_i0_reset),
    .io_d(AsyncResetRegVec_w1_i0_io_d),
    .io_q(AsyncResetRegVec_w1_i0_io_q),
    .io_en(AsyncResetRegVec_w1_i0_io_en)
  );
  assign _T = io_deq_ready & io_deq_valid; 
  assign source_ready = AsyncValidSync_2_io_out; 
  assign _T_1 = source_ready == 1'h0; 
  assign _GEN_8 = {{3'd0}, _T}; 
  assign _T_4 = ridx_bin_io_q + _GEN_8; 
  assign _T_5 = _T_1 ? 4'h0 : _T_4; 
  assign _T_6 = _T_5[3:1]; 
  assign _GEN_9 = {{1'd0}, _T_6}; 
  assign ridx = _T_5 ^ _GEN_9; 
  assign widx = widx_gray_io_q; 
  assign _T_7 = ridx != widx; 
  assign valid = source_ready & _T_7; 
  assign _T_8 = ridx[2:0]; 
  assign _T_9 = ridx[3]; 
  assign _T_10 = {_T_9, 2'h0}; 
  assign index = _T_8 ^ _T_10; 
  assign _GEN_1 = 3'h1 == index ? io_async_mem_1 : io_async_mem_0; 
  assign _GEN_2 = 3'h2 == index ? io_async_mem_2 : _GEN_1; 
  assign _GEN_3 = 3'h3 == index ? io_async_mem_3 : _GEN_2; 
  assign _GEN_4 = 3'h4 == index ? io_async_mem_4 : _GEN_3; 
  assign _GEN_5 = 3'h5 == index ? io_async_mem_5 : _GEN_4; 
  assign _GEN_6 = 3'h6 == index ? io_async_mem_6 : _GEN_5; 
  assign _GEN_7 = 3'h7 == index ? io_async_mem_7 : _GEN_6; 
  assign valid_reg_1 = valid_reg_io_q; 
  assign _T_14 = io_async_safe_source_reset_n == 1'h0; 
  assign io_deq_valid = valid_reg_1 & source_ready; 
  assign io_deq_bits = deq_bits_reg_io_q; 
  assign io_async_ridx = ridx_gray_io_q; 
  assign io_async_safe_ridx_valid = AsyncValidSync_io_out; 
  assign io_async_safe_sink_reset_n = reset == 1'h0; 
  assign ridx_bin_clock = clock; 
  assign ridx_bin_reset = reset; 
  assign ridx_bin_io_d = _T_1 ? 4'h0 : _T_4; 
  assign ridx_bin_io_en = 1'h1; 
  assign widx_gray_clock = clock; 
  assign widx_gray_reset = reset; 
  assign widx_gray_io_d = io_async_widx; 
  assign deq_bits_reg_clock = clock; 
  assign deq_bits_reg_io_d = valid ? _GEN_7 : io_deq_bits; 
  assign valid_reg_clock = clock; 
  assign valid_reg_reset = reset; 
  assign valid_reg_io_d = source_ready & _T_7; 
  assign valid_reg_io_en = 1'h1; 
  assign ridx_gray_clock = clock; 
  assign ridx_gray_reset = reset; 
  assign ridx_gray_io_d = _T_5 ^ _GEN_9; 
  assign ridx_gray_io_en = 1'h1; 
  assign AsyncValidSync_clock = clock; 
  assign AsyncValidSync_reset = reset | _T_14; 
  assign AsyncValidSync_io_in = 1'h1; 
  assign AsyncValidSync_1_clock = clock; 
  assign AsyncValidSync_1_reset = reset | _T_14; 
  assign AsyncValidSync_1_io_in = io_async_safe_widx_valid; 
  assign AsyncValidSync_2_clock = clock; 
  assign AsyncValidSync_2_reset = reset; 
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out; 
  assign AsyncResetRegVec_w1_i0_clock = clock; 
  assign AsyncResetRegVec_w1_i0_reset = reset; 
  assign AsyncResetRegVec_w1_i0_io_d = io_async_widx == io_async_ridx; 
  assign AsyncResetRegVec_w1_i0_io_en = 1'h1; 
endmodule
module dual_AsyncQueueSource_5( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [19:0] io_enq_bits_a, 
  input  [19:0] io_enq_bits_b, 
  input  [19:0] io_enq_bits_c, 
  input  [19:0] io_enq_bits_d, 
  input  [19:0] io_enq_bits_e, 
  output [19:0] io_async_mem_0_a, 
  output [19:0] io_async_mem_0_b, 
  output [19:0] io_async_mem_0_c, 
  output [19:0] io_async_mem_0_d, 
  output [19:0] io_async_mem_0_e, 
  input         io_async_ridx, 
  output        io_async_widx, 
  input         io_async_safe_ridx_valid, 
  output        io_async_safe_widx_valid, 
  output        io_async_safe_source_reset_n, 
  input         io_async_safe_sink_reset_n 
);
  wire  widx_bin_clock; 
  wire  widx_bin_reset; 
  wire  widx_bin_io_d; 
  wire  widx_bin_io_q; 
  wire  widx_bin_io_en; 
  wire  ridx_gray_clock; 
  wire  ridx_gray_reset; 
  wire  ridx_gray_io_d; 
  wire  ridx_gray_io_q; 
  wire  ready_reg_clock; 
  wire  ready_reg_reset; 
  wire  ready_reg_io_d; 
  wire  ready_reg_io_q; 
  wire  ready_reg_io_en; 
  wire  widx_gray_clock; 
  wire  widx_gray_reset; 
  wire  widx_gray_io_d; 
  wire  widx_gray_io_q; 
  wire  widx_gray_io_en; 
  wire  AsyncValidSync_clock; 
  wire  AsyncValidSync_reset; 
  wire  AsyncValidSync_io_in; 
  wire  AsyncValidSync_io_out; 
  wire  AsyncValidSync_1_clock; 
  wire  AsyncValidSync_1_reset; 
  wire  AsyncValidSync_1_io_in; 
  wire  AsyncValidSync_1_io_out; 
  wire  AsyncValidSync_2_clock; 
  wire  AsyncValidSync_2_reset; 
  wire  AsyncValidSync_2_io_in; 
  wire  AsyncValidSync_2_io_out; 
  reg [19:0] mem_0_a; 
  reg [31:0] _RAND_0;
  reg [19:0] mem_0_b; 
  reg [31:0] _RAND_1;
  reg [19:0] mem_0_c; 
  reg [31:0] _RAND_2;
  reg [19:0] mem_0_d; 
  reg [31:0] _RAND_3;
  reg [19:0] mem_0_e; 
  reg [31:0] _RAND_4;
  wire  _T; 
  wire  sink_ready; 
  wire  _T_1; 
  wire  _T_4; 
  wire  widx; 
  wire  ridx; 
  wire  _T_7; 
  wire  _T_8; 
  wire  ready_reg_1; 
  wire  _T_12; 
  dual_AsyncResetRegVec_w1_i0 widx_bin ( 
    .clock(widx_bin_clock),
    .reset(widx_bin_reset),
    .io_d(widx_bin_io_d),
    .io_q(widx_bin_io_q),
    .io_en(widx_bin_io_en)
  );
  dual_AsyncResetSynchronizerShiftReg_w1_d3_i0 ridx_gray ( 
    .clock(ridx_gray_clock),
    .reset(ridx_gray_reset),
    .io_d(ridx_gray_io_d),
    .io_q(ridx_gray_io_q)
  );
  dual_AsyncResetRegVec_w1_i0 ready_reg ( 
    .clock(ready_reg_clock),
    .reset(ready_reg_reset),
    .io_d(ready_reg_io_d),
    .io_q(ready_reg_io_q),
    .io_en(ready_reg_io_en)
  );
  dual_AsyncResetRegVec_w1_i0 widx_gray ( 
    .clock(widx_gray_clock),
    .reset(widx_gray_reset),
    .io_d(widx_gray_io_d),
    .io_q(widx_gray_io_q),
    .io_en(widx_gray_io_en)
  );
  dual_AsyncValidSync AsyncValidSync ( 
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_in(AsyncValidSync_io_in),
    .io_out(AsyncValidSync_io_out)
  );
  dual_AsyncValidSync_1 AsyncValidSync_1 ( 
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  dual_AsyncValidSync_2 AsyncValidSync_2 ( 
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  assign _T = io_enq_ready & io_enq_valid; 
  assign sink_ready = AsyncValidSync_2_io_out; 
  assign _T_1 = sink_ready == 1'h0; 
  assign _T_4 = widx_bin_io_q + _T; 
  assign widx = _T_1 ? 1'h0 : _T_4; 
  assign ridx = ridx_gray_io_q; 
  assign _T_7 = ridx ^ 1'h1; 
  assign _T_8 = widx != _T_7; 
  assign ready_reg_1 = ready_reg_io_q; 
  assign _T_12 = io_async_safe_sink_reset_n == 1'h0; 
  assign io_enq_ready = ready_reg_1 & sink_ready; 
  assign io_async_mem_0_a = mem_0_a; 
  assign io_async_mem_0_b = mem_0_b; 
  assign io_async_mem_0_c = mem_0_c; 
  assign io_async_mem_0_d = mem_0_d; 
  assign io_async_mem_0_e = mem_0_e; 
  assign io_async_widx = widx_gray_io_q; 
  assign io_async_safe_widx_valid = AsyncValidSync_io_out; 
  assign io_async_safe_source_reset_n = reset == 1'h0; 
  assign widx_bin_clock = clock; 
  assign widx_bin_reset = reset; 
  assign widx_bin_io_d = _T_1 ? 1'h0 : _T_4; 
  assign widx_bin_io_en = 1'h1; 
  assign ridx_gray_clock = clock; 
  assign ridx_gray_reset = reset; 
  assign ridx_gray_io_d = io_async_ridx; 
  assign ready_reg_clock = clock; 
  assign ready_reg_reset = reset; 
  assign ready_reg_io_d = sink_ready & _T_8; 
  assign ready_reg_io_en = 1'h1; 
  assign widx_gray_clock = clock; 
  assign widx_gray_reset = reset; 
  assign widx_gray_io_d = _T_1 ? 1'h0 : _T_4; 
  assign widx_gray_io_en = 1'h1; 
  assign AsyncValidSync_clock = clock; 
  assign AsyncValidSync_reset = reset | _T_12; 
  assign AsyncValidSync_io_in = 1'h1; 
  assign AsyncValidSync_1_clock = clock; 
  assign AsyncValidSync_1_reset = reset | _T_12; 
  assign AsyncValidSync_1_io_in = io_async_safe_ridx_valid; 
  assign AsyncValidSync_2_clock = clock; 
  assign AsyncValidSync_2_reset = reset; 
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0_a = _RAND_0[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_0_b = _RAND_1[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_0_c = _RAND_2[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_0_d = _RAND_3[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  mem_0_e = _RAND_4[19:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (_T) begin
      mem_0_a <= io_enq_bits_a;
    end
    if (_T) begin
      mem_0_b <= io_enq_bits_b;
    end
    if (_T) begin
      mem_0_c <= io_enq_bits_c;
    end
    if (_T) begin
      mem_0_d <= io_enq_bits_d;
    end
    if (_T) begin
      mem_0_e <= io_enq_bits_e;
    end
  end
endmodule
module dual_AsyncQueueSource( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [31:0] io_enq_bits, 
  output [31:0] io_async_mem_0, 
  output [31:0] io_async_mem_1, 
  output [31:0] io_async_mem_2, 
  output [31:0] io_async_mem_3, 
  output [31:0] io_async_mem_4, 
  output [31:0] io_async_mem_5, 
  output [31:0] io_async_mem_6, 
  output [31:0] io_async_mem_7, 
  input  [3:0]  io_async_ridx, 
  output [3:0]  io_async_widx, 
  input         io_async_safe_ridx_valid, 
  output        io_async_safe_widx_valid, 
  output        io_async_safe_source_reset_n, 
  input         io_async_safe_sink_reset_n 
);
  wire  widx_bin_clock; 
  wire  widx_bin_reset; 
  wire [3:0] widx_bin_io_d; 
  wire [3:0] widx_bin_io_q; 
  wire  widx_bin_io_en; 
  wire  ridx_gray_clock; 
  wire  ridx_gray_reset; 
  wire [3:0] ridx_gray_io_d; 
  wire [3:0] ridx_gray_io_q; 
  wire  ready_reg_clock; 
  wire  ready_reg_reset; 
  wire  ready_reg_io_d; 
  wire  ready_reg_io_q; 
  wire  ready_reg_io_en; 
  wire  widx_gray_clock; 
  wire  widx_gray_reset; 
  wire [3:0] widx_gray_io_d; 
  wire [3:0] widx_gray_io_q; 
  wire  widx_gray_io_en; 
  wire  AsyncValidSync_clock; 
  wire  AsyncValidSync_reset; 
  wire  AsyncValidSync_io_in; 
  wire  AsyncValidSync_io_out; 
  wire  AsyncValidSync_1_clock; 
  wire  AsyncValidSync_1_reset; 
  wire  AsyncValidSync_1_io_in; 
  wire  AsyncValidSync_1_io_out; 
  wire  AsyncValidSync_2_clock; 
  wire  AsyncValidSync_2_reset; 
  wire  AsyncValidSync_2_io_in; 
  wire  AsyncValidSync_2_io_out; 
  reg [31:0] mem_0; 
  reg [31:0] _RAND_0;
  reg [31:0] mem_1; 
  reg [31:0] _RAND_1;
  reg [31:0] mem_2; 
  reg [31:0] _RAND_2;
  reg [31:0] mem_3; 
  reg [31:0] _RAND_3;
  reg [31:0] mem_4; 
  reg [31:0] _RAND_4;
  reg [31:0] mem_5; 
  reg [31:0] _RAND_5;
  reg [31:0] mem_6; 
  reg [31:0] _RAND_6;
  reg [31:0] mem_7; 
  reg [31:0] _RAND_7;
  wire  _T; 
  wire  sink_ready; 
  wire  _T_1; 
  wire [3:0] _GEN_16; 
  wire [3:0] _T_4; 
  wire [3:0] _T_5; 
  wire [2:0] _T_6; 
  wire [3:0] _GEN_17; 
  wire [3:0] widx; 
  wire [3:0] ridx; 
  wire [3:0] _T_7; 
  wire  _T_8; 
  wire [2:0] _T_9; 
  wire  _T_10; 
  wire [2:0] _T_11; 
  wire [2:0] index; 
  wire  ready_reg_1; 
  wire  _T_15; 
  dual_AsyncResetRegVec_w4_i0 widx_bin ( 
    .clock(widx_bin_clock),
    .reset(widx_bin_reset),
    .io_d(widx_bin_io_d),
    .io_q(widx_bin_io_q),
    .io_en(widx_bin_io_en)
  );
  dual_AsyncResetSynchronizerShiftReg_w4_d3_i0 ridx_gray ( 
    .clock(ridx_gray_clock),
    .reset(ridx_gray_reset),
    .io_d(ridx_gray_io_d),
    .io_q(ridx_gray_io_q)
  );
  dual_AsyncResetRegVec_w1_i0 ready_reg ( 
    .clock(ready_reg_clock),
    .reset(ready_reg_reset),
    .io_d(ready_reg_io_d),
    .io_q(ready_reg_io_q),
    .io_en(ready_reg_io_en)
  );
  dual_AsyncResetRegVec_w4_i0 widx_gray ( 
    .clock(widx_gray_clock),
    .reset(widx_gray_reset),
    .io_d(widx_gray_io_d),
    .io_q(widx_gray_io_q),
    .io_en(widx_gray_io_en)
  );
  dual_AsyncValidSync AsyncValidSync ( 
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_in(AsyncValidSync_io_in),
    .io_out(AsyncValidSync_io_out)
  );
  dual_AsyncValidSync_1 AsyncValidSync_1 ( 
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  dual_AsyncValidSync_2 AsyncValidSync_2 ( 
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  assign _T = io_enq_ready & io_enq_valid; 
  assign sink_ready = AsyncValidSync_2_io_out; 
  assign _T_1 = sink_ready == 1'h0; 
  assign _GEN_16 = {{3'd0}, _T}; 
  assign _T_4 = widx_bin_io_q + _GEN_16; 
  assign _T_5 = _T_1 ? 4'h0 : _T_4; 
  assign _T_6 = _T_5[3:1]; 
  assign _GEN_17 = {{1'd0}, _T_6}; 
  assign widx = _T_5 ^ _GEN_17; 
  assign ridx = ridx_gray_io_q; 
  assign _T_7 = ridx ^ 4'hc; 
  assign _T_8 = widx != _T_7; 
  assign _T_9 = io_async_widx[2:0]; 
  assign _T_10 = io_async_widx[3]; 
  assign _T_11 = {_T_10, 2'h0}; 
  assign index = _T_9 ^ _T_11; 
  assign ready_reg_1 = ready_reg_io_q; 
  assign _T_15 = io_async_safe_sink_reset_n == 1'h0; 
  assign io_enq_ready = ready_reg_1 & sink_ready; 
  assign io_async_mem_0 = mem_0; 
  assign io_async_mem_1 = mem_1; 
  assign io_async_mem_2 = mem_2; 
  assign io_async_mem_3 = mem_3; 
  assign io_async_mem_4 = mem_4; 
  assign io_async_mem_5 = mem_5; 
  assign io_async_mem_6 = mem_6; 
  assign io_async_mem_7 = mem_7; 
  assign io_async_widx = widx_gray_io_q; 
  assign io_async_safe_widx_valid = AsyncValidSync_io_out; 
  assign io_async_safe_source_reset_n = reset == 1'h0; 
  assign widx_bin_clock = clock; 
  assign widx_bin_reset = reset; 
  assign widx_bin_io_d = _T_1 ? 4'h0 : _T_4; 
  assign widx_bin_io_en = 1'h1; 
  assign ridx_gray_clock = clock; 
  assign ridx_gray_reset = reset; 
  assign ridx_gray_io_d = io_async_ridx; 
  assign ready_reg_clock = clock; 
  assign ready_reg_reset = reset; 
  assign ready_reg_io_d = sink_ready & _T_8; 
  assign ready_reg_io_en = 1'h1; 
  assign widx_gray_clock = clock; 
  assign widx_gray_reset = reset; 
  assign widx_gray_io_d = _T_5 ^ _GEN_17; 
  assign widx_gray_io_en = 1'h1; 
  assign AsyncValidSync_clock = clock; 
  assign AsyncValidSync_reset = reset | _T_15; 
  assign AsyncValidSync_io_in = 1'h1; 
  assign AsyncValidSync_1_clock = clock; 
  assign AsyncValidSync_1_reset = reset | _T_15; 
  assign AsyncValidSync_1_io_in = io_async_safe_ridx_valid; 
  assign AsyncValidSync_2_clock = clock; 
  assign AsyncValidSync_2_reset = reset; 
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  mem_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  mem_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mem_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mem_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (_T) begin
      if (3'h0 == index) begin
        mem_0 <= io_enq_bits;
      end
    end
    if (_T) begin
      if (3'h1 == index) begin
        mem_1 <= io_enq_bits;
      end
    end
    if (_T) begin
      if (3'h2 == index) begin
        mem_2 <= io_enq_bits;
      end
    end
    if (_T) begin
      if (3'h3 == index) begin
        mem_3 <= io_enq_bits;
      end
    end
    if (_T) begin
      if (3'h4 == index) begin
        mem_4 <= io_enq_bits;
      end
    end
    if (_T) begin
      if (3'h5 == index) begin
        mem_5 <= io_enq_bits;
      end
    end
    if (_T) begin
      if (3'h6 == index) begin
        mem_6 <= io_enq_bits;
      end
    end
    if (_T) begin
      if (3'h7 == index) begin
        mem_7 <= io_enq_bits;
      end
    end
  end
endmodule
module dual_AsyncResetReg (d, q, en, clk, rst);
parameter RESET_VALUE = 0;

input  wire d;
output reg  q;
input  wire en;
input  wire clk;
input  wire rst;

   // There is a lot of initialization
   // here you don't normally find in Verilog
   // async registers because of scenarios in which reset
   // is not actually asserted cleanly at time 0,
   // and we want to make sure to properly model
   // that, yet Chisel codebase is absolutely intolerant
   // of Xs.
`ifndef SYNTHESIS
  initial begin:B0
    `ifdef RANDOMIZE
    integer    initvar;
    reg [31:0] _RAND;
    _RAND = {1{$random}};
    q = _RAND[0];
    `endif // RANDOMIZE
    if (rst) begin
      q = RESET_VALUE;
    end 
  end
`endif

   always @(posedge clk or posedge rst) begin

      if (rst) begin
         q <= RESET_VALUE;
      end else if (en) begin
         q <= d;
      end
   end
 
endmodule // dual_AsyncResetReg

/* verilator lint_off UNOPTFLAT */

module dual_AsyncResetRegVec_w1_i0( 
  input   clock, 
  input   reset, 
  input   io_d, 
  output  io_q, 
  input   io_en 
);
  wire  reg_0_d; 
  wire  reg_0_q; 
  wire  reg_0_en; 
  wire  reg_0_clk; 
  wire  reg_0_rst; 
  dual_AsyncResetReg #(.RESET_VALUE(0)) reg_0 ( 
    .d(reg_0_d),
    .q(reg_0_q),
    .en(reg_0_en),
    .clk(reg_0_clk),
    .rst(reg_0_rst)
  );
  assign io_q = reg_0_q; 
  assign reg_0_d = io_d; 
  assign reg_0_en = io_en; 
  assign reg_0_clk = clock; 
  assign reg_0_rst = reset; 
endmodule
module dual_AsyncResetRegVec_w4_i0( 
  input        clock, 
  input        reset, 
  input  [3:0] io_d, 
  output [3:0] io_q, 
  input        io_en 
);
  wire  reg_0_d; 
  wire  reg_0_q; 
  wire  reg_0_en; 
  wire  reg_0_clk; 
  wire  reg_0_rst; 
  wire  reg_1_d; 
  wire  reg_1_q; 
  wire  reg_1_en; 
  wire  reg_1_clk; 
  wire  reg_1_rst; 
  wire  reg_2_d; 
  wire  reg_2_q; 
  wire  reg_2_en; 
  wire  reg_2_clk; 
  wire  reg_2_rst; 
  wire  reg_3_d; 
  wire  reg_3_q; 
  wire  reg_3_en; 
  wire  reg_3_clk; 
  wire  reg_3_rst; 
  wire [1:0] _T_4; 
  wire [1:0] _T_5; 
  dual_AsyncResetReg #(.RESET_VALUE(0)) reg_0 ( 
    .d(reg_0_d),
    .q(reg_0_q),
    .en(reg_0_en),
    .clk(reg_0_clk),
    .rst(reg_0_rst)
  );
  dual_AsyncResetReg #(.RESET_VALUE(0)) reg_1 ( 
    .d(reg_1_d),
    .q(reg_1_q),
    .en(reg_1_en),
    .clk(reg_1_clk),
    .rst(reg_1_rst)
  );
  dual_AsyncResetReg #(.RESET_VALUE(0)) reg_2 ( 
    .d(reg_2_d),
    .q(reg_2_q),
    .en(reg_2_en),
    .clk(reg_2_clk),
    .rst(reg_2_rst)
  );
  dual_AsyncResetReg #(.RESET_VALUE(0)) reg_3 ( 
    .d(reg_3_d),
    .q(reg_3_q),
    .en(reg_3_en),
    .clk(reg_3_clk),
    .rst(reg_3_rst)
  );
  assign _T_4 = {reg_1_q,reg_0_q}; 
  assign _T_5 = {reg_3_q,reg_2_q}; 
  assign io_q = {_T_5,_T_4}; 
  assign reg_0_d = io_d[0]; 
  assign reg_0_en = io_en; 
  assign reg_0_clk = clock; 
  assign reg_0_rst = reset; 
  assign reg_1_d = io_d[1]; 
  assign reg_1_en = io_en; 
  assign reg_1_clk = clock; 
  assign reg_1_rst = reset; 
  assign reg_2_d = io_d[2]; 
  assign reg_2_en = io_en; 
  assign reg_2_clk = clock; 
  assign reg_2_rst = reset; 
  assign reg_3_d = io_d[3]; 
  assign reg_3_en = io_en; 
  assign reg_3_clk = clock; 
  assign reg_3_rst = reset; 
endmodule
module dual_AsyncResetSynchronizerShiftReg_w1_d1_i0( 
  input   clock, 
  input   reset, 
  input   io_d, 
  output  io_q 
);
  wire  sync_0_clock; 
  wire  sync_0_reset; 
  wire  sync_0_io_d; 
  wire  sync_0_io_q; 
  wire  sync_0_io_en; 
  dual_AsyncResetRegVec_w1_i0 sync_0 ( 
    .clock(sync_0_clock),
    .reset(sync_0_reset),
    .io_d(sync_0_io_d),
    .io_q(sync_0_io_q),
    .io_en(sync_0_io_en)
  );
  assign io_q = sync_0_io_q; 
  assign sync_0_clock = clock; 
  assign sync_0_reset = reset; 
  assign sync_0_io_d = io_d; 
  assign sync_0_io_en = 1'h1; 
endmodule
module dual_AsyncResetSynchronizerShiftReg_w1_d3_i0( 
  input   clock, 
  input   reset, 
  input   io_d, 
  output  io_q 
);
  wire  sync_0_clock; 
  wire  sync_0_reset; 
  wire  sync_0_io_d; 
  wire  sync_0_io_q; 
  wire  sync_0_io_en; 
  wire  sync_1_clock; 
  wire  sync_1_reset; 
  wire  sync_1_io_d; 
  wire  sync_1_io_q; 
  wire  sync_1_io_en; 
  wire  sync_2_clock; 
  wire  sync_2_reset; 
  wire  sync_2_io_d; 
  wire  sync_2_io_q; 
  wire  sync_2_io_en; 
  dual_AsyncResetRegVec_w1_i0 sync_0 ( 
    .clock(sync_0_clock),
    .reset(sync_0_reset),
    .io_d(sync_0_io_d),
    .io_q(sync_0_io_q),
    .io_en(sync_0_io_en)
  );
  dual_AsyncResetRegVec_w1_i0 sync_1 ( 
    .clock(sync_1_clock),
    .reset(sync_1_reset),
    .io_d(sync_1_io_d),
    .io_q(sync_1_io_q),
    .io_en(sync_1_io_en)
  );
  dual_AsyncResetRegVec_w1_i0 sync_2 ( 
    .clock(sync_2_clock),
    .reset(sync_2_reset),
    .io_d(sync_2_io_d),
    .io_q(sync_2_io_q),
    .io_en(sync_2_io_en)
  );
  assign io_q = sync_0_io_q; 
  assign sync_0_clock = clock; 
  assign sync_0_reset = reset; 
  assign sync_0_io_d = sync_1_io_q; 
  assign sync_0_io_en = 1'h1; 
  assign sync_1_clock = clock; 
  assign sync_1_reset = reset; 
  assign sync_1_io_d = sync_2_io_q; 
  assign sync_1_io_en = 1'h1; 
  assign sync_2_clock = clock; 
  assign sync_2_reset = reset; 
  assign sync_2_io_d = io_d; 
  assign sync_2_io_en = 1'h1; 
endmodule
module dual_AsyncResetSynchronizerShiftReg_w1_d4_i0( 
  input   clock, 
  input   reset, 
  input   io_d, 
  output  io_q 
);
  wire  sync_0_clock; 
  wire  sync_0_reset; 
  wire  sync_0_io_d; 
  wire  sync_0_io_q; 
  wire  sync_0_io_en; 
  wire  sync_1_clock; 
  wire  sync_1_reset; 
  wire  sync_1_io_d; 
  wire  sync_1_io_q; 
  wire  sync_1_io_en; 
  wire  sync_2_clock; 
  wire  sync_2_reset; 
  wire  sync_2_io_d; 
  wire  sync_2_io_q; 
  wire  sync_2_io_en; 
  wire  sync_3_clock; 
  wire  sync_3_reset; 
  wire  sync_3_io_d; 
  wire  sync_3_io_q; 
  wire  sync_3_io_en; 
  dual_AsyncResetRegVec_w1_i0 sync_0 ( 
    .clock(sync_0_clock),
    .reset(sync_0_reset),
    .io_d(sync_0_io_d),
    .io_q(sync_0_io_q),
    .io_en(sync_0_io_en)
  );
  dual_AsyncResetRegVec_w1_i0 sync_1 ( 
    .clock(sync_1_clock),
    .reset(sync_1_reset),
    .io_d(sync_1_io_d),
    .io_q(sync_1_io_q),
    .io_en(sync_1_io_en)
  );
  dual_AsyncResetRegVec_w1_i0 sync_2 ( 
    .clock(sync_2_clock),
    .reset(sync_2_reset),
    .io_d(sync_2_io_d),
    .io_q(sync_2_io_q),
    .io_en(sync_2_io_en)
  );
  dual_AsyncResetRegVec_w1_i0 sync_3 ( 
    .clock(sync_3_clock),
    .reset(sync_3_reset),
    .io_d(sync_3_io_d),
    .io_q(sync_3_io_q),
    .io_en(sync_3_io_en)
  );
  assign io_q = sync_0_io_q; 
  assign sync_0_clock = clock; 
  assign sync_0_reset = reset; 
  assign sync_0_io_d = sync_1_io_q; 
  assign sync_0_io_en = 1'h1; 
  assign sync_1_clock = clock; 
  assign sync_1_reset = reset; 
  assign sync_1_io_d = sync_2_io_q; 
  assign sync_1_io_en = 1'h1; 
  assign sync_2_clock = clock; 
  assign sync_2_reset = reset; 
  assign sync_2_io_d = sync_3_io_q; 
  assign sync_2_io_en = 1'h1; 
  assign sync_3_clock = clock; 
  assign sync_3_reset = reset; 
  assign sync_3_io_d = io_d; 
  assign sync_3_io_en = 1'h1; 
endmodule
module dual_AsyncResetSynchronizerShiftReg_w4_d3_i0( 
  input        clock, 
  input        reset, 
  input  [3:0] io_d, 
  output [3:0] io_q 
);
  wire  sync_0_clock; 
  wire  sync_0_reset; 
  wire [3:0] sync_0_io_d; 
  wire [3:0] sync_0_io_q; 
  wire  sync_0_io_en; 
  wire  sync_1_clock; 
  wire  sync_1_reset; 
  wire [3:0] sync_1_io_d; 
  wire [3:0] sync_1_io_q; 
  wire  sync_1_io_en; 
  wire  sync_2_clock; 
  wire  sync_2_reset; 
  wire [3:0] sync_2_io_d; 
  wire [3:0] sync_2_io_q; 
  wire  sync_2_io_en; 
  dual_AsyncResetRegVec_w4_i0 sync_0 ( 
    .clock(sync_0_clock),
    .reset(sync_0_reset),
    .io_d(sync_0_io_d),
    .io_q(sync_0_io_q),
    .io_en(sync_0_io_en)
  );
  dual_AsyncResetRegVec_w4_i0 sync_1 ( 
    .clock(sync_1_clock),
    .reset(sync_1_reset),
    .io_d(sync_1_io_d),
    .io_q(sync_1_io_q),
    .io_en(sync_1_io_en)
  );
  dual_AsyncResetRegVec_w4_i0 sync_2 ( 
    .clock(sync_2_clock),
    .reset(sync_2_reset),
    .io_d(sync_2_io_d),
    .io_q(sync_2_io_q),
    .io_en(sync_2_io_en)
  );
  assign io_q = sync_0_io_q; 
  assign sync_0_clock = clock; 
  assign sync_0_reset = reset; 
  assign sync_0_io_d = sync_1_io_q; 
  assign sync_0_io_en = 1'h1; 
  assign sync_1_clock = clock; 
  assign sync_1_reset = reset; 
  assign sync_1_io_d = sync_2_io_q; 
  assign sync_1_io_en = 1'h1; 
  assign sync_2_clock = clock; 
  assign sync_2_reset = reset; 
  assign sync_2_io_d = io_d; 
  assign sync_2_io_en = 1'h1; 
endmodule
module dual_AsyncValidSync_1( 
  input   clock, 
  input   reset, 
  input   io_in, 
  output  io_out 
);
  wire  sink_extend_clock; 
  wire  sink_extend_reset; 
  wire  sink_extend_io_d; 
  wire  sink_extend_io_q; 
  dual_AsyncResetSynchronizerShiftReg_w1_d1_i0 sink_extend ( 
    .clock(sink_extend_clock),
    .reset(sink_extend_reset),
    .io_d(sink_extend_io_d),
    .io_q(sink_extend_io_q)
  );
  assign io_out = sink_extend_io_q; 
  assign sink_extend_clock = clock; 
  assign sink_extend_reset = reset; 
  assign sink_extend_io_d = io_in; 
endmodule
module dual_AsyncValidSync_2( 
  input   clock, 
  input   reset, 
  input   io_in, 
  output  io_out 
);
  wire  sink_valid_clock; 
  wire  sink_valid_reset; 
  wire  sink_valid_io_d; 
  wire  sink_valid_io_q; 
  dual_AsyncResetSynchronizerShiftReg_w1_d3_i0 sink_valid ( 
    .clock(sink_valid_clock),
    .reset(sink_valid_reset),
    .io_d(sink_valid_io_d),
    .io_q(sink_valid_io_q)
  );
  assign io_out = sink_valid_io_q; 
  assign sink_valid_clock = clock; 
  assign sink_valid_reset = reset; 
  assign sink_valid_io_d = io_in; 
endmodule
module dual_AsyncValidSync( 
  input   clock, 
  input   reset, 
  input   io_in, 
  output  io_out 
);
  wire  source_valid_clock; 
  wire  source_valid_reset; 
  wire  source_valid_io_d; 
  wire  source_valid_io_q; 
  dual_AsyncResetSynchronizerShiftReg_w1_d4_i0 source_valid ( 
    .clock(source_valid_clock),
    .reset(source_valid_reset),
    .io_d(source_valid_io_d),
    .io_q(source_valid_io_q)
  );
  assign io_out = source_valid_io_q; 
  assign source_valid_clock = clock; 
  assign source_valid_reset = reset; 
  assign source_valid_io_d = io_in; 
endmodule
module dual_AXI4Buffer( 
  input         clock, 
  input         reset, 
  output        auto_in_awready, 
  input         auto_in_awvalid, 
  input  [30:0] auto_in_awaddr, 
  input  [7:0]  auto_in_awlen, 
  input  [2:0]  auto_in_awsize, 
  input  [1:0]  auto_in_awburst, 
  input         auto_in_awlock, 
  input  [3:0]  auto_in_awcache, 
  input  [2:0]  auto_in_awprot, 
  input  [3:0]  auto_in_awqos, 
  input  [63:0] auto_in_awinstret, 
  output        auto_in_wready, 
  input         auto_in_wvalid, 
  input  [63:0] auto_in_wdata, 
  input  [7:0]  auto_in_wstrb, 
  input         auto_in_wlast, 
  input         auto_in_bready, 
  output        auto_in_bvalid, 
  output [1:0]  auto_in_bresp, 
  output        auto_in_arready, 
  input         auto_in_arvalid, 
  input  [30:0] auto_in_araddr, 
  input  [7:0]  auto_in_arlen, 
  input  [2:0]  auto_in_arsize, 
  input  [1:0]  auto_in_arburst, 
  input         auto_in_arlock, 
  input  [3:0]  auto_in_arcache, 
  input  [2:0]  auto_in_arprot, 
  input  [3:0]  auto_in_arqos, 
  input  [63:0] auto_in_arinstret, 
  input         auto_in_rready, 
  output        auto_in_rvalid, 
  output [63:0] auto_in_rdata, 
  output [1:0]  auto_in_rresp, 
  output        auto_in_rlast, 
  input         auto_out_awready, 
  output        auto_out_awvalid, 
  output        auto_out_awid, 
  output [30:0] auto_out_awaddr, 
  output [7:0]  auto_out_awlen, 
  output [2:0]  auto_out_awsize, 
  output [1:0]  auto_out_awburst, 
  output        auto_out_awlock, 
  output [3:0]  auto_out_awcache, 
  output [2:0]  auto_out_awprot, 
  output [3:0]  auto_out_awqos, 
  output [63:0] auto_out_awinstret, 
  input         auto_out_wready, 
  output        auto_out_wvalid, 
  output [63:0] auto_out_wdata, 
  output [7:0]  auto_out_wstrb, 
  output        auto_out_wlast, 
  output        auto_out_bready, 
  input         auto_out_bvalid, 
  input  [1:0]  auto_out_bresp, 
  input         auto_out_arready, 
  output        auto_out_arvalid, 
  output        auto_out_arid, 
  output [30:0] auto_out_araddr, 
  output [7:0]  auto_out_arlen, 
  output [2:0]  auto_out_arsize, 
  output [1:0]  auto_out_arburst, 
  output        auto_out_arlock, 
  output [3:0]  auto_out_arcache, 
  output [2:0]  auto_out_arprot, 
  output [3:0]  auto_out_arqos, 
  output [63:0] auto_out_arinstret, 
  output        auto_out_rready, 
  input         auto_out_rvalid, 
  input  [63:0] auto_out_rdata, 
  input  [1:0]  auto_out_rresp, 
  input         auto_out_rlast 
);
  wire  Queue_clock; 
  wire  Queue_reset; 
  wire  Queue_io_enq_ready; 
  wire  Queue_io_enq_valid; 
  wire [30:0] Queue_io_enq_bits_addr; 
  wire [7:0] Queue_io_enq_bits_len; 
  wire [2:0] Queue_io_enq_bits_size; 
  wire [1:0] Queue_io_enq_bits_burst; 
  wire  Queue_io_enq_bits_lock; 
  wire [3:0] Queue_io_enq_bits_cache; 
  wire [2:0] Queue_io_enq_bits_prot; 
  wire [3:0] Queue_io_enq_bits_qos; 
  wire [63:0] Queue_io_enq_bits_instret; 
  wire  Queue_io_deq_ready; 
  wire  Queue_io_deq_valid; 
  wire  Queue_io_deq_bits_id; 
  wire [30:0] Queue_io_deq_bits_addr; 
  wire [7:0] Queue_io_deq_bits_len; 
  wire [2:0] Queue_io_deq_bits_size; 
  wire [1:0] Queue_io_deq_bits_burst; 
  wire  Queue_io_deq_bits_lock; 
  wire [3:0] Queue_io_deq_bits_cache; 
  wire [2:0] Queue_io_deq_bits_prot; 
  wire [3:0] Queue_io_deq_bits_qos; 
  wire [63:0] Queue_io_deq_bits_instret; 
  wire  Queue_1_clock; 
  wire  Queue_1_reset; 
  wire  Queue_1_io_enq_ready; 
  wire  Queue_1_io_enq_valid; 
  wire [63:0] Queue_1_io_enq_bits_data; 
  wire [7:0] Queue_1_io_enq_bits_strb; 
  wire  Queue_1_io_enq_bits_last; 
  wire  Queue_1_io_deq_ready; 
  wire  Queue_1_io_deq_valid; 
  wire [63:0] Queue_1_io_deq_bits_data; 
  wire [7:0] Queue_1_io_deq_bits_strb; 
  wire  Queue_1_io_deq_bits_last; 
  wire  Queue_2_clock; 
  wire  Queue_2_reset; 
  wire  Queue_2_io_enq_ready; 
  wire  Queue_2_io_enq_valid; 
  wire [1:0] Queue_2_io_enq_bits_resp; 
  wire  Queue_2_io_deq_ready; 
  wire  Queue_2_io_deq_valid; 
  wire [1:0] Queue_2_io_deq_bits_resp; 
  wire  Queue_3_clock; 
  wire  Queue_3_reset; 
  wire  Queue_3_io_enq_ready; 
  wire  Queue_3_io_enq_valid; 
  wire [30:0] Queue_3_io_enq_bits_addr; 
  wire [7:0] Queue_3_io_enq_bits_len; 
  wire [2:0] Queue_3_io_enq_bits_size; 
  wire [1:0] Queue_3_io_enq_bits_burst; 
  wire  Queue_3_io_enq_bits_lock; 
  wire [3:0] Queue_3_io_enq_bits_cache; 
  wire [2:0] Queue_3_io_enq_bits_prot; 
  wire [3:0] Queue_3_io_enq_bits_qos; 
  wire [63:0] Queue_3_io_enq_bits_instret; 
  wire  Queue_3_io_deq_ready; 
  wire  Queue_3_io_deq_valid; 
  wire  Queue_3_io_deq_bits_id; 
  wire [30:0] Queue_3_io_deq_bits_addr; 
  wire [7:0] Queue_3_io_deq_bits_len; 
  wire [2:0] Queue_3_io_deq_bits_size; 
  wire [1:0] Queue_3_io_deq_bits_burst; 
  wire  Queue_3_io_deq_bits_lock; 
  wire [3:0] Queue_3_io_deq_bits_cache; 
  wire [2:0] Queue_3_io_deq_bits_prot; 
  wire [3:0] Queue_3_io_deq_bits_qos; 
  wire [63:0] Queue_3_io_deq_bits_instret; 
  wire  Queue_4_clock; 
  wire  Queue_4_reset; 
  wire  Queue_4_io_enq_ready; 
  wire  Queue_4_io_enq_valid; 
  wire [63:0] Queue_4_io_enq_bits_data; 
  wire [1:0] Queue_4_io_enq_bits_resp; 
  wire  Queue_4_io_enq_bits_last; 
  wire  Queue_4_io_deq_ready; 
  wire  Queue_4_io_deq_valid; 
  wire [63:0] Queue_4_io_deq_bits_data; 
  wire [1:0] Queue_4_io_deq_bits_resp; 
  wire  Queue_4_io_deq_bits_last; 
  dual_Queue_48 dual_Queue ( 
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_addr(Queue_io_enq_bits_addr),
    .io_enq_bits_len(Queue_io_enq_bits_len),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_burst(Queue_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_io_enq_bits_qos),
    .io_enq_bits_instret(Queue_io_enq_bits_instret),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_addr(Queue_io_deq_bits_addr),
    .io_deq_bits_len(Queue_io_deq_bits_len),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_burst(Queue_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_io_deq_bits_qos),
    .io_deq_bits_instret(Queue_io_deq_bits_instret)
  );
  dual_Queue_49 Queue_1 ( 
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_strb(Queue_1_io_enq_bits_strb),
    .io_enq_bits_last(Queue_1_io_enq_bits_last),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_strb(Queue_1_io_deq_bits_strb),
    .io_deq_bits_last(Queue_1_io_deq_bits_last)
  );
  dual_Queue_50 dual_Queue_2 ( 
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_resp(Queue_2_io_enq_bits_resp),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_resp(Queue_2_io_deq_bits_resp)
  );
  dual_Queue_48 Queue_3 ( 
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_addr(Queue_3_io_enq_bits_addr),
    .io_enq_bits_len(Queue_3_io_enq_bits_len),
    .io_enq_bits_size(Queue_3_io_enq_bits_size),
    .io_enq_bits_burst(Queue_3_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_3_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_3_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_3_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_3_io_enq_bits_qos),
    .io_enq_bits_instret(Queue_3_io_enq_bits_instret),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_id(Queue_3_io_deq_bits_id),
    .io_deq_bits_addr(Queue_3_io_deq_bits_addr),
    .io_deq_bits_len(Queue_3_io_deq_bits_len),
    .io_deq_bits_size(Queue_3_io_deq_bits_size),
    .io_deq_bits_burst(Queue_3_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_3_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_3_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_3_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_3_io_deq_bits_qos),
    .io_deq_bits_instret(Queue_3_io_deq_bits_instret)
  );
  dual_Queue_52 dual_Queue_4 ( 
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_data(Queue_4_io_enq_bits_data),
    .io_enq_bits_resp(Queue_4_io_enq_bits_resp),
    .io_enq_bits_last(Queue_4_io_enq_bits_last),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_data(Queue_4_io_deq_bits_data),
    .io_deq_bits_resp(Queue_4_io_deq_bits_resp),
    .io_deq_bits_last(Queue_4_io_deq_bits_last)
  );
  assign auto_in_awready = Queue_io_enq_ready; 
  assign auto_in_wready = Queue_1_io_enq_ready; 
  assign auto_in_bvalid = Queue_2_io_deq_valid; 
  assign auto_in_bresp = Queue_2_io_deq_bits_resp; 
  assign auto_in_arready = Queue_3_io_enq_ready; 
  assign auto_in_rvalid = Queue_4_io_deq_valid; 
  assign auto_in_rdata = Queue_4_io_deq_bits_data; 
  assign auto_in_rresp = Queue_4_io_deq_bits_resp; 
  assign auto_in_rlast = Queue_4_io_deq_bits_last; 
  assign auto_out_awvalid = Queue_io_deq_valid; 
  assign auto_out_awid = Queue_io_deq_bits_id; 
  assign auto_out_awaddr = Queue_io_deq_bits_addr; 
  assign auto_out_awlen = Queue_io_deq_bits_len; 
  assign auto_out_awsize = Queue_io_deq_bits_size; 
  assign auto_out_awburst = Queue_io_deq_bits_burst; 
  assign auto_out_awlock = Queue_io_deq_bits_lock; 
  assign auto_out_awcache = Queue_io_deq_bits_cache; 
  assign auto_out_awprot = Queue_io_deq_bits_prot; 
  assign auto_out_awqos = Queue_io_deq_bits_qos; 
  assign auto_out_awinstret = Queue_io_deq_bits_instret; 
  assign auto_out_wvalid = Queue_1_io_deq_valid; 
  assign auto_out_wdata = Queue_1_io_deq_bits_data; 
  assign auto_out_wstrb = Queue_1_io_deq_bits_strb; 
  assign auto_out_wlast = Queue_1_io_deq_bits_last; 
  assign auto_out_bready = Queue_2_io_enq_ready; 
  assign auto_out_arvalid = Queue_3_io_deq_valid; 
  assign auto_out_arid = Queue_3_io_deq_bits_id; 
  assign auto_out_araddr = Queue_3_io_deq_bits_addr; 
  assign auto_out_arlen = Queue_3_io_deq_bits_len; 
  assign auto_out_arsize = Queue_3_io_deq_bits_size; 
  assign auto_out_arburst = Queue_3_io_deq_bits_burst; 
  assign auto_out_arlock = Queue_3_io_deq_bits_lock; 
  assign auto_out_arcache = Queue_3_io_deq_bits_cache; 
  assign auto_out_arprot = Queue_3_io_deq_bits_prot; 
  assign auto_out_arqos = Queue_3_io_deq_bits_qos; 
  assign auto_out_arinstret = Queue_3_io_deq_bits_instret; 
  assign auto_out_rready = Queue_4_io_enq_ready; 
  assign Queue_clock = clock; 
  assign Queue_reset = reset; 
  assign Queue_io_enq_valid = auto_in_awvalid; 
  assign Queue_io_enq_bits_addr = auto_in_awaddr; 
  assign Queue_io_enq_bits_len = auto_in_awlen; 
  assign Queue_io_enq_bits_size = auto_in_awsize; 
  assign Queue_io_enq_bits_burst = auto_in_awburst; 
  assign Queue_io_enq_bits_lock = auto_in_awlock; 
  assign Queue_io_enq_bits_cache = auto_in_awcache; 
  assign Queue_io_enq_bits_prot = auto_in_awprot; 
  assign Queue_io_enq_bits_qos = auto_in_awqos; 
  assign Queue_io_enq_bits_instret = auto_in_awinstret; 
  assign Queue_io_deq_ready = auto_out_awready; 
  assign Queue_1_clock = clock; 
  assign Queue_1_reset = reset; 
  assign Queue_1_io_enq_valid = auto_in_wvalid; 
  assign Queue_1_io_enq_bits_data = auto_in_wdata; 
  assign Queue_1_io_enq_bits_strb = auto_in_wstrb; 
  assign Queue_1_io_enq_bits_last = auto_in_wlast; 
  assign Queue_1_io_deq_ready = auto_out_wready; 
  assign Queue_2_clock = clock; 
  assign Queue_2_reset = reset; 
  assign Queue_2_io_enq_valid = auto_out_bvalid; 
  assign Queue_2_io_enq_bits_resp = auto_out_bresp; 
  assign Queue_2_io_deq_ready = auto_in_bready; 
  assign Queue_3_clock = clock; 
  assign Queue_3_reset = reset; 
  assign Queue_3_io_enq_valid = auto_in_arvalid; 
  assign Queue_3_io_enq_bits_addr = auto_in_araddr; 
  assign Queue_3_io_enq_bits_len = auto_in_arlen; 
  assign Queue_3_io_enq_bits_size = auto_in_arsize; 
  assign Queue_3_io_enq_bits_burst = auto_in_arburst; 
  assign Queue_3_io_enq_bits_lock = auto_in_arlock; 
  assign Queue_3_io_enq_bits_cache = auto_in_arcache; 
  assign Queue_3_io_enq_bits_prot = auto_in_arprot; 
  assign Queue_3_io_enq_bits_qos = auto_in_arqos; 
  assign Queue_3_io_enq_bits_instret = auto_in_arinstret; 
  assign Queue_3_io_deq_ready = auto_out_arready; 
  assign Queue_4_clock = clock; 
  assign Queue_4_reset = reset; 
  assign Queue_4_io_enq_valid = auto_out_rvalid; 
  assign Queue_4_io_enq_bits_data = auto_out_rdata; 
  assign Queue_4_io_enq_bits_resp = auto_out_rresp; 
  assign Queue_4_io_enq_bits_last = auto_out_rlast; 
  assign Queue_4_io_deq_ready = auto_in_rready; 
endmodule
module dual_AXI4Deinterleaver( 
  input         clock, 
  input         reset, 
  output        auto_in_awready, 
  input         auto_in_awvalid, 
  input  [30:0] auto_in_awaddr, 
  input  [7:0]  auto_in_awlen, 
  input  [2:0]  auto_in_awsize, 
  input  [1:0]  auto_in_awburst, 
  input         auto_in_awlock, 
  input  [3:0]  auto_in_awcache, 
  input  [2:0]  auto_in_awprot, 
  input  [3:0]  auto_in_awqos, 
  input  [15:0] auto_in_awuser, 
  input  [63:0] auto_in_awinstret, 
  output        auto_in_wready, 
  input         auto_in_wvalid, 
  input  [63:0] auto_in_wdata, 
  input  [7:0]  auto_in_wstrb, 
  input         auto_in_wlast, 
  input         auto_in_bready, 
  output        auto_in_bvalid, 
  output [1:0]  auto_in_bresp, 
  output [15:0] auto_in_buser, 
  output        auto_in_arready, 
  input         auto_in_arvalid, 
  input  [30:0] auto_in_araddr, 
  input  [7:0]  auto_in_arlen, 
  input  [2:0]  auto_in_arsize, 
  input  [1:0]  auto_in_arburst, 
  input         auto_in_arlock, 
  input  [3:0]  auto_in_arcache, 
  input  [2:0]  auto_in_arprot, 
  input  [3:0]  auto_in_arqos, 
  input  [15:0] auto_in_aruser, 
  input  [63:0] auto_in_arinstret, 
  input         auto_in_rready, 
  output        auto_in_rvalid, 
  output [63:0] auto_in_rdata, 
  output [1:0]  auto_in_rresp, 
  output [15:0] auto_in_ruser, 
  output        auto_in_rlast, 
  input         auto_out_awready, 
  output        auto_out_awvalid, 
  output [30:0] auto_out_awaddr, 
  output [7:0]  auto_out_awlen, 
  output [2:0]  auto_out_awsize, 
  output [1:0]  auto_out_awburst, 
  output        auto_out_awlock, 
  output [3:0]  auto_out_awcache, 
  output [2:0]  auto_out_awprot, 
  output [3:0]  auto_out_awqos, 
  output [15:0] auto_out_awuser, 
  output [63:0] auto_out_awinstret, 
  input         auto_out_wready, 
  output        auto_out_wvalid, 
  output [63:0] auto_out_wdata, 
  output [7:0]  auto_out_wstrb, 
  output        auto_out_wlast, 
  output        auto_out_bready, 
  input         auto_out_bvalid, 
  input  [1:0]  auto_out_bresp, 
  input  [15:0] auto_out_buser, 
  input         auto_out_arready, 
  output        auto_out_arvalid, 
  output [30:0] auto_out_araddr, 
  output [7:0]  auto_out_arlen, 
  output [2:0]  auto_out_arsize, 
  output [1:0]  auto_out_arburst, 
  output        auto_out_arlock, 
  output [3:0]  auto_out_arcache, 
  output [2:0]  auto_out_arprot, 
  output [3:0]  auto_out_arqos, 
  output [15:0] auto_out_aruser, 
  output [63:0] auto_out_arinstret, 
  output        auto_out_rready, 
  input         auto_out_rvalid, 
  input  [63:0] auto_out_rdata, 
  input  [1:0]  auto_out_rresp, 
  input  [15:0] auto_out_ruser, 
  input         auto_out_rlast 
);
  wire  Queue_clock; 
  wire  Queue_reset; 
  wire  Queue_io_enq_ready; 
  wire  Queue_io_enq_valid; 
  wire [63:0] Queue_io_enq_bits_data; 
  wire [1:0] Queue_io_enq_bits_resp; 
  wire [15:0] Queue_io_enq_bits_user; 
  wire  Queue_io_enq_bits_last; 
  wire  Queue_io_deq_ready; 
  wire  Queue_io_deq_valid; 
  wire [63:0] Queue_io_deq_bits_data; 
  wire [1:0] Queue_io_deq_bits_resp; 
  wire [15:0] Queue_io_deq_bits_user; 
  wire  Queue_io_deq_bits_last; 
  reg  _T_2; 
  reg [31:0] _RAND_0;
  reg [3:0] _T_4; 
  reg [31:0] _RAND_1;
  wire  _T_42_0; 
  wire  _T_6; 
  wire  _T_8; 
  wire  _T_9; 
  wire  _T_39_0_last; 
  wire  _T_11; 
  wire [3:0] _GEN_2; 
  wire [3:0] _T_13; 
  wire [3:0] _GEN_3; 
  wire [3:0] _T_15; 
  wire  _T_16; 
  wire  _T_17; 
  wire  _T_18; 
  wire  _T_20; 
  wire  _T_21; 
  wire  _T_22; 
  wire  _T_23; 
  wire  _T_24; 
  wire  _T_26; 
  wire  _T_27; 
  wire  _T_28; 
  wire  _T_33; 
  wire  _T_36; 
  dual_Queue_55 dual_Queue ( 
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_resp(Queue_io_enq_bits_resp),
    .io_enq_bits_user(Queue_io_enq_bits_user),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_resp(Queue_io_deq_bits_resp),
    .io_deq_bits_user(Queue_io_deq_bits_user),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign _T_42_0 = Queue_io_enq_ready; 
  assign _T_6 = _T_42_0 & auto_out_rvalid; 
  assign _T_8 = _T_6 & auto_out_rlast; 
  assign _T_9 = auto_in_rready & _T_2; 
  assign _T_39_0_last = Queue_io_deq_bits_last; 
  assign _T_11 = _T_9 & _T_39_0_last; 
  assign _GEN_2 = {{3'd0}, _T_8}; 
  assign _T_13 = _T_4 + _GEN_2; 
  assign _GEN_3 = {{3'd0}, _T_11}; 
  assign _T_15 = _T_13 - _GEN_3; 
  assign _T_16 = _T_11 == 1'h0; 
  assign _T_17 = _T_4 != 4'h0; 
  assign _T_18 = _T_16 | _T_17; 
  assign _T_20 = _T_18 | reset; 
  assign _T_21 = _T_20 == 1'h0; 
  assign _T_22 = _T_8 == 1'h0; 
  assign _T_23 = _T_4 != 4'h8; 
  assign _T_24 = _T_22 | _T_23; 
  assign _T_26 = _T_24 | reset; 
  assign _T_27 = _T_26 == 1'h0; 
  assign _T_28 = _T_15 != 4'h0; 
  assign _T_33 = _T_2 == 1'h0; 
  assign _T_36 = _T_33 | _T_11; 
  assign auto_in_awready = auto_out_awready; 
  assign auto_in_wready = auto_out_wready; 
  assign auto_in_bvalid = auto_out_bvalid; 
  assign auto_in_bresp = auto_out_bresp; 
  assign auto_in_buser = auto_out_buser; 
  assign auto_in_arready = auto_out_arready; 
  assign auto_in_rvalid = _T_2; 
  assign auto_in_rdata = Queue_io_deq_bits_data; 
  assign auto_in_rresp = Queue_io_deq_bits_resp; 
  assign auto_in_ruser = Queue_io_deq_bits_user; 
  assign auto_in_rlast = Queue_io_deq_bits_last; 
  assign auto_out_awvalid = auto_in_awvalid; 
  assign auto_out_awaddr = auto_in_awaddr; 
  assign auto_out_awlen = auto_in_awlen; 
  assign auto_out_awsize = auto_in_awsize; 
  assign auto_out_awburst = auto_in_awburst; 
  assign auto_out_awlock = auto_in_awlock; 
  assign auto_out_awcache = auto_in_awcache; 
  assign auto_out_awprot = auto_in_awprot; 
  assign auto_out_awqos = auto_in_awqos; 
  assign auto_out_awuser = auto_in_awuser; 
  assign auto_out_awinstret = auto_in_awinstret; 
  assign auto_out_wvalid = auto_in_wvalid; 
  assign auto_out_wdata = auto_in_wdata; 
  assign auto_out_wstrb = auto_in_wstrb; 
  assign auto_out_wlast = auto_in_wlast; 
  assign auto_out_bready = auto_in_bready; 
  assign auto_out_arvalid = auto_in_arvalid; 
  assign auto_out_araddr = auto_in_araddr; 
  assign auto_out_arlen = auto_in_arlen; 
  assign auto_out_arsize = auto_in_arsize; 
  assign auto_out_arburst = auto_in_arburst; 
  assign auto_out_arlock = auto_in_arlock; 
  assign auto_out_arcache = auto_in_arcache; 
  assign auto_out_arprot = auto_in_arprot; 
  assign auto_out_arqos = auto_in_arqos; 
  assign auto_out_aruser = auto_in_aruser; 
  assign auto_out_arinstret = auto_in_arinstret; 
  assign auto_out_rready = Queue_io_enq_ready; 
  assign Queue_clock = clock; 
  assign Queue_reset = reset; 
  assign Queue_io_enq_valid = auto_out_rvalid; 
  assign Queue_io_enq_bits_data = auto_out_rdata; 
  assign Queue_io_enq_bits_resp = auto_out_rresp; 
  assign Queue_io_enq_bits_user = auto_out_ruser; 
  assign Queue_io_enq_bits_last = auto_out_rlast; 
  assign Queue_io_deq_ready = auto_in_rready & _T_2; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_4 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_2 <= 1'h0;
    end else begin
      if (_T_36) begin
        _T_2 <= _T_28;
      end
    end
    if (reset) begin
      _T_4 <= 4'h0;
    end else begin
      _T_4 <= _T_15;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:69 assert (!dec || count =/= UInt(0))\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_21) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_27) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:70 assert (!inc || count =/= UInt(beats))\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_27) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_AXI4Fragmenter( 
  input         clock, 
  input         reset, 
  output        auto_in_awready, 
  input         auto_in_awvalid, 
  input         auto_in_awid, 
  input  [31:0] auto_in_awaddr, 
  input  [7:0]  auto_in_awlen, 
  input  [2:0]  auto_in_awsize, 
  input  [1:0]  auto_in_awburst, 
  input  [15:0] auto_in_awuser, 
  output        auto_in_wready, 
  input         auto_in_wvalid, 
  input  [63:0] auto_in_wdata, 
  input  [7:0]  auto_in_wstrb, 
  input         auto_in_wlast, 
  input         auto_in_bready, 
  output        auto_in_bvalid, 
  output        auto_in_bid, 
  output [1:0]  auto_in_bresp, 
  output [15:0] auto_in_buser, 
  output        auto_in_arready, 
  input         auto_in_arvalid, 
  input         auto_in_arid, 
  input  [31:0] auto_in_araddr, 
  input  [7:0]  auto_in_arlen, 
  input  [2:0]  auto_in_arsize, 
  input  [1:0]  auto_in_arburst, 
  input  [15:0] auto_in_aruser, 
  input         auto_in_rready, 
  output        auto_in_rvalid, 
  output        auto_in_rid, 
  output [63:0] auto_in_rdata, 
  output [1:0]  auto_in_rresp, 
  output [15:0] auto_in_ruser, 
  output        auto_in_rlast, 
  input         auto_out_awready, 
  output        auto_out_awvalid, 
  output        auto_out_awid, 
  output [31:0] auto_out_awaddr, 
  output [7:0]  auto_out_awlen, 
  output [2:0]  auto_out_awsize, 
  output [16:0] auto_out_awuser, 
  input         auto_out_wready, 
  output        auto_out_wvalid, 
  output [63:0] auto_out_wdata, 
  output [7:0]  auto_out_wstrb, 
  output        auto_out_wlast, 
  output        auto_out_bready, 
  input         auto_out_bvalid, 
  input         auto_out_bid, 
  input  [1:0]  auto_out_bresp, 
  input  [16:0] auto_out_buser, 
  input         auto_out_arready, 
  output        auto_out_arvalid, 
  output        auto_out_arid, 
  output [31:0] auto_out_araddr, 
  output [7:0]  auto_out_arlen, 
  output [2:0]  auto_out_arsize, 
  output [16:0] auto_out_aruser, 
  output        auto_out_rready, 
  input         auto_out_rvalid, 
  input         auto_out_rid, 
  input  [63:0] auto_out_rdata, 
  input  [1:0]  auto_out_rresp, 
  input  [16:0] auto_out_ruser, 
  input         auto_out_rlast 
);
  wire  Queue_clock; 
  wire  Queue_reset; 
  wire  Queue_io_enq_ready; 
  wire  Queue_io_enq_valid; 
  wire  Queue_io_enq_bits_id; 
  wire [31:0] Queue_io_enq_bits_addr; 
  wire [7:0] Queue_io_enq_bits_len; 
  wire [2:0] Queue_io_enq_bits_size; 
  wire [1:0] Queue_io_enq_bits_burst; 
  wire [15:0] Queue_io_enq_bits_user; 
  wire  Queue_io_deq_ready; 
  wire  Queue_io_deq_valid; 
  wire  Queue_io_deq_bits_id; 
  wire [31:0] Queue_io_deq_bits_addr; 
  wire [7:0] Queue_io_deq_bits_len; 
  wire [2:0] Queue_io_deq_bits_size; 
  wire [1:0] Queue_io_deq_bits_burst; 
  wire [15:0] Queue_io_deq_bits_user; 
  wire  Queue_1_clock; 
  wire  Queue_1_reset; 
  wire  Queue_1_io_enq_ready; 
  wire  Queue_1_io_enq_valid; 
  wire  Queue_1_io_enq_bits_id; 
  wire [31:0] Queue_1_io_enq_bits_addr; 
  wire [7:0] Queue_1_io_enq_bits_len; 
  wire [2:0] Queue_1_io_enq_bits_size; 
  wire [1:0] Queue_1_io_enq_bits_burst; 
  wire [15:0] Queue_1_io_enq_bits_user; 
  wire  Queue_1_io_deq_ready; 
  wire  Queue_1_io_deq_valid; 
  wire  Queue_1_io_deq_bits_id; 
  wire [31:0] Queue_1_io_deq_bits_addr; 
  wire [7:0] Queue_1_io_deq_bits_len; 
  wire [2:0] Queue_1_io_deq_bits_size; 
  wire [1:0] Queue_1_io_deq_bits_burst; 
  wire [15:0] Queue_1_io_deq_bits_user; 
  wire  Queue_2_clock; 
  wire  Queue_2_reset; 
  wire  Queue_2_io_enq_ready; 
  wire  Queue_2_io_enq_valid; 
  wire [63:0] Queue_2_io_enq_bits_data; 
  wire [7:0] Queue_2_io_enq_bits_strb; 
  wire  Queue_2_io_enq_bits_last; 
  wire  Queue_2_io_deq_ready; 
  wire  Queue_2_io_deq_valid; 
  wire [63:0] Queue_2_io_deq_bits_data; 
  wire [7:0] Queue_2_io_deq_bits_strb; 
  wire  Queue_2_io_deq_bits_last; 
  reg  _T_4; 
  reg [31:0] _RAND_0;
  reg [31:0] _T_5; 
  reg [31:0] _RAND_1;
  reg [7:0] _T_6; 
  reg [31:0] _RAND_2;
  wire [7:0] _T_2_bits_len; 
  wire [7:0] _T_7; 
  wire [31:0] _T_2_bits_addr; 
  wire [31:0] _T_8; 
  wire [7:0] _T_10; 
  wire [6:0] _T_16; 
  wire [7:0] _GEN_16; 
  wire [7:0] _T_17; 
  wire [5:0] _T_18; 
  wire [7:0] _GEN_17; 
  wire [7:0] _T_19; 
  wire [3:0] _T_20; 
  wire [7:0] _GEN_18; 
  wire [7:0] _T_21; 
  wire [6:0] _T_23; 
  wire [7:0] _T_24; 
  wire [8:0] _T_25; 
  wire [7:0] _T_26; 
  wire [7:0] _T_27; 
  wire [9:0] _T_28; 
  wire [7:0] _T_29; 
  wire [7:0] _T_30; 
  wire [11:0] _T_31; 
  wire [7:0] _T_32; 
  wire [7:0] _T_33; 
  wire [7:0] _T_35; 
  wire [7:0] _GEN_19; 
  wire [7:0] _T_36; 
  wire [8:0] _T_37; 
  wire [7:0] _T_38; 
  wire [7:0] _T_39; 
  wire [9:0] _T_40; 
  wire [7:0] _T_41; 
  wire [7:0] _T_42; 
  wire [11:0] _T_43; 
  wire [7:0] _T_44; 
  wire [7:0] _T_45; 
  wire [7:0] _T_47; 
  wire [7:0] _T_48; 
  wire [7:0] _T_49; 
  wire [1:0] _T_2_bits_burst; 
  wire  _T_50; 
  wire [2:0] _T_2_bits_size; 
  wire  _T_51; 
  wire  _T_52; 
  wire [7:0] _T_53; 
  wire [8:0] _T_54; 
  wire [8:0] _T_55; 
  wire [8:0] _T_56; 
  wire [8:0] _T_57; 
  wire [8:0] _T_58; 
  wire [15:0] _GEN_20; 
  wire [15:0] _T_59; 
  wire [31:0] _GEN_21; 
  wire [31:0] _T_61; 
  wire [15:0] _T_62; 
  wire [22:0] _GEN_22; 
  wire [22:0] _T_63; 
  wire [14:0] _T_64; 
  wire  _T_66; 
  wire [31:0] _GEN_23; 
  wire [31:0] _T_67; 
  wire [31:0] _T_68; 
  wire [31:0] _T_69; 
  wire [31:0] _T_70; 
  wire [31:0] _T_71; 
  wire  _T_73; 
  wire [31:0] _T_75; 
  wire [9:0] _T_77; 
  wire [2:0] _T_78; 
  wire [2:0] _T_79; 
  wire [31:0] _GEN_25; 
  wire [31:0] _T_80; 
  wire  _T_2_valid; 
  wire  _T_82; 
  wire  _T_83; 
  wire [8:0] _GEN_26; 
  wire [8:0] _T_85; 
  wire [8:0] _GEN_4; 
  reg  _T_88; 
  reg [31:0] _RAND_3;
  reg [31:0] _T_89; 
  reg [31:0] _RAND_4;
  reg [7:0] _T_90; 
  reg [31:0] _RAND_5;
  wire [7:0] _T_86_bits_len; 
  wire [7:0] _T_91; 
  wire [31:0] _T_86_bits_addr; 
  wire [31:0] _T_92; 
  wire [7:0] _T_94; 
  wire [6:0] _T_100; 
  wire [7:0] _GEN_27; 
  wire [7:0] _T_101; 
  wire [5:0] _T_102; 
  wire [7:0] _GEN_28; 
  wire [7:0] _T_103; 
  wire [3:0] _T_104; 
  wire [7:0] _GEN_29; 
  wire [7:0] _T_105; 
  wire [6:0] _T_107; 
  wire [7:0] _T_108; 
  wire [8:0] _T_109; 
  wire [7:0] _T_110; 
  wire [7:0] _T_111; 
  wire [9:0] _T_112; 
  wire [7:0] _T_113; 
  wire [7:0] _T_114; 
  wire [11:0] _T_115; 
  wire [7:0] _T_116; 
  wire [7:0] _T_117; 
  wire [7:0] _T_119; 
  wire [7:0] _GEN_30; 
  wire [7:0] _T_120; 
  wire [8:0] _T_121; 
  wire [7:0] _T_122; 
  wire [7:0] _T_123; 
  wire [9:0] _T_124; 
  wire [7:0] _T_125; 
  wire [7:0] _T_126; 
  wire [11:0] _T_127; 
  wire [7:0] _T_128; 
  wire [7:0] _T_129; 
  wire [7:0] _T_131; 
  wire [7:0] _T_132; 
  wire [7:0] _T_133; 
  wire [1:0] _T_86_bits_burst; 
  wire  _T_134; 
  wire [2:0] _T_86_bits_size; 
  wire  _T_135; 
  wire  _T_136; 
  wire [7:0] _T_137; 
  wire [8:0] _T_138; 
  wire [8:0] _T_139; 
  wire [8:0] _T_140; 
  wire [8:0] _T_141; 
  wire [8:0] _T_142; 
  wire [15:0] _GEN_31; 
  wire [15:0] _T_143; 
  wire [31:0] _GEN_32; 
  wire [31:0] _T_145; 
  wire [15:0] _T_146; 
  wire [22:0] _GEN_33; 
  wire [22:0] _T_147; 
  wire [14:0] _T_148; 
  wire  _T_150; 
  wire [31:0] _GEN_34; 
  wire [31:0] _T_151; 
  wire [31:0] _T_152; 
  wire [31:0] _T_153; 
  wire [31:0] _T_154; 
  wire [31:0] _T_155; 
  wire  _T_157; 
  reg [8:0] _T_184; 
  reg [31:0] _RAND_6;
  wire  _T_185; 
  reg  _T_172; 
  reg [31:0] _RAND_7;
  wire  _T_179; 
  wire  _T_180; 
  wire [31:0] _T_159; 
  wire [9:0] _T_161; 
  wire [2:0] _T_162; 
  wire [2:0] _T_163; 
  wire [31:0] _GEN_36; 
  wire [31:0] _T_164; 
  wire  _T_86_valid; 
  wire  _T_166; 
  wire  _T_167; 
  wire [8:0] _GEN_37; 
  wire [8:0] _T_169; 
  wire [8:0] _GEN_9; 
  wire [15:0] _T_2_bits_user; 
  wire  _T_181; 
  wire  _T_182; 
  wire  _T_175; 
  wire  _T_178; 
  wire  _T_176; 
  wire [15:0] _T_86_bits_user; 
  wire [8:0] _T_186; 
  wire [8:0] _T_187; 
  wire  _T_188; 
  wire  _T_170_valid; 
  wire  _T_199; 
  wire  _T_200; 
  wire  _T_201; 
  wire  _T_189; 
  wire [8:0] _GEN_38; 
  wire [8:0] _T_191; 
  wire  _T_193; 
  wire  _T_194; 
  wire  _T_195; 
  wire  _T_197; 
  wire  _T_198; 
  wire  _T_205; 
  wire  _T_170_bits_last; 
  wire  _T_206; 
  wire  _T_207; 
  wire  _T_208; 
  wire  _T_210; 
  wire  _T_211; 
  wire  _T_212; 
  wire  _T_215; 
  wire  _T_217; 
  wire  _T_218; 
  reg [1:0] _T_221_0; 
  reg [31:0] _RAND_8;
  reg [1:0] _T_221_1; 
  reg [31:0] _RAND_9;
  wire [1:0] _GEN_13; 
  wire [1:0] _T_224; 
  wire  _T_226; 
  wire  _T_227; 
  wire  _T_228; 
  wire  _T_229; 
  wire [1:0] _T_230; 
  wire  _T_233; 
  wire [1:0] _T_234; 
  dual_Queue_64 dual_Queue ( 
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_addr(Queue_io_enq_bits_addr),
    .io_enq_bits_len(Queue_io_enq_bits_len),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_burst(Queue_io_enq_bits_burst),
    .io_enq_bits_user(Queue_io_enq_bits_user),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_addr(Queue_io_deq_bits_addr),
    .io_deq_bits_len(Queue_io_deq_bits_len),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_burst(Queue_io_deq_bits_burst),
    .io_deq_bits_user(Queue_io_deq_bits_user)
  );
  dual_Queue_64 Queue_1 ( 
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_id(Queue_1_io_enq_bits_id),
    .io_enq_bits_addr(Queue_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_burst(Queue_1_io_enq_bits_burst),
    .io_enq_bits_user(Queue_1_io_enq_bits_user),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_id(Queue_1_io_deq_bits_id),
    .io_deq_bits_addr(Queue_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_1_io_deq_bits_burst),
    .io_deq_bits_user(Queue_1_io_deq_bits_user)
  );
  dual_Queue_46 dual_Queue_2 ( 
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_data(Queue_2_io_enq_bits_data),
    .io_enq_bits_strb(Queue_2_io_enq_bits_strb),
    .io_enq_bits_last(Queue_2_io_enq_bits_last),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_data(Queue_2_io_deq_bits_data),
    .io_deq_bits_strb(Queue_2_io_deq_bits_strb),
    .io_deq_bits_last(Queue_2_io_deq_bits_last)
  );
  assign _T_2_bits_len = Queue_io_deq_bits_len; 
  assign _T_7 = _T_4 ? _T_6 : _T_2_bits_len; 
  assign _T_2_bits_addr = Queue_io_deq_bits_addr; 
  assign _T_8 = _T_4 ? _T_5 : _T_2_bits_addr; 
  assign _T_10 = _T_8[10:3]; 
  assign _T_16 = _T_7[7:1]; 
  assign _GEN_16 = {{1'd0}, _T_16}; 
  assign _T_17 = _T_7 | _GEN_16; 
  assign _T_18 = _T_17[7:2]; 
  assign _GEN_17 = {{2'd0}, _T_18}; 
  assign _T_19 = _T_17 | _GEN_17; 
  assign _T_20 = _T_19[7:4]; 
  assign _GEN_18 = {{4'd0}, _T_20}; 
  assign _T_21 = _T_19 | _GEN_18; 
  assign _T_23 = _T_21[7:1]; 
  assign _T_24 = ~ _T_7; 
  assign _T_25 = {_T_24, 1'h0}; 
  assign _T_26 = _T_25[7:0]; 
  assign _T_27 = _T_24 | _T_26; 
  assign _T_28 = {_T_27, 2'h0}; 
  assign _T_29 = _T_28[7:0]; 
  assign _T_30 = _T_27 | _T_29; 
  assign _T_31 = {_T_30, 4'h0}; 
  assign _T_32 = _T_31[7:0]; 
  assign _T_33 = _T_30 | _T_32; 
  assign _T_35 = ~ _T_33; 
  assign _GEN_19 = {{1'd0}, _T_23}; 
  assign _T_36 = _GEN_19 | _T_35; 
  assign _T_37 = {_T_10, 1'h0}; 
  assign _T_38 = _T_37[7:0]; 
  assign _T_39 = _T_10 | _T_38; 
  assign _T_40 = {_T_39, 2'h0}; 
  assign _T_41 = _T_40[7:0]; 
  assign _T_42 = _T_39 | _T_41; 
  assign _T_43 = {_T_42, 4'h0}; 
  assign _T_44 = _T_43[7:0]; 
  assign _T_45 = _T_42 | _T_44; 
  assign _T_47 = ~ _T_45; 
  assign _T_48 = _T_36 & _T_47; 
  assign _T_49 = _T_48 & 8'h7; 
  assign _T_2_bits_burst = Queue_io_deq_bits_burst; 
  assign _T_50 = _T_2_bits_burst == 2'h0; 
  assign _T_2_bits_size = Queue_io_deq_bits_size; 
  assign _T_51 = _T_2_bits_size != 3'h3; 
  assign _T_52 = _T_50 | _T_51; 
  assign _T_53 = _T_52 ? 8'h0 : _T_49; 
  assign _T_54 = {_T_53, 1'h0}; 
  assign _T_55 = _T_54 | 9'h1; 
  assign _T_56 = {1'h0,_T_53}; 
  assign _T_57 = ~ _T_56; 
  assign _T_58 = _T_55 & _T_57; 
  assign _GEN_20 = {{7'd0}, _T_58}; 
  assign _T_59 = _GEN_20 << _T_2_bits_size; 
  assign _GEN_21 = {{16'd0}, _T_59}; 
  assign _T_61 = _T_8 + _GEN_21; 
  assign _T_62 = {_T_2_bits_len,8'hff}; 
  assign _GEN_22 = {{7'd0}, _T_62}; 
  assign _T_63 = _GEN_22 << _T_2_bits_size; 
  assign _T_64 = _T_63[22:8]; 
  assign _T_66 = _T_2_bits_burst == 2'h2; 
  assign _GEN_23 = {{17'd0}, _T_64}; 
  assign _T_67 = _T_61 & _GEN_23; 
  assign _T_68 = ~ _T_2_bits_addr; 
  assign _T_69 = _T_68 | _GEN_23; 
  assign _T_70 = ~ _T_69; 
  assign _T_71 = _T_67 | _T_70; 
  assign _T_73 = _T_53 == _T_7; 
  assign _T_75 = ~ _T_8; 
  assign _T_77 = 10'h7 << _T_2_bits_size; 
  assign _T_78 = _T_77[2:0]; 
  assign _T_79 = ~ _T_78; 
  assign _GEN_25 = {{29'd0}, _T_79}; 
  assign _T_80 = _T_75 | _GEN_25; 
  assign _T_2_valid = Queue_io_deq_valid; 
  assign _T_82 = auto_out_arready & _T_2_valid; 
  assign _T_83 = _T_73 == 1'h0; 
  assign _GEN_26 = {{1'd0}, _T_7}; 
  assign _T_85 = _GEN_26 - _T_58; 
  assign _GEN_4 = _T_82 ? _T_85 : {{1'd0}, _T_6}; 
  assign _T_86_bits_len = Queue_1_io_deq_bits_len; 
  assign _T_91 = _T_88 ? _T_90 : _T_86_bits_len; 
  assign _T_86_bits_addr = Queue_1_io_deq_bits_addr; 
  assign _T_92 = _T_88 ? _T_89 : _T_86_bits_addr; 
  assign _T_94 = _T_92[10:3]; 
  assign _T_100 = _T_91[7:1]; 
  assign _GEN_27 = {{1'd0}, _T_100}; 
  assign _T_101 = _T_91 | _GEN_27; 
  assign _T_102 = _T_101[7:2]; 
  assign _GEN_28 = {{2'd0}, _T_102}; 
  assign _T_103 = _T_101 | _GEN_28; 
  assign _T_104 = _T_103[7:4]; 
  assign _GEN_29 = {{4'd0}, _T_104}; 
  assign _T_105 = _T_103 | _GEN_29; 
  assign _T_107 = _T_105[7:1]; 
  assign _T_108 = ~ _T_91; 
  assign _T_109 = {_T_108, 1'h0}; 
  assign _T_110 = _T_109[7:0]; 
  assign _T_111 = _T_108 | _T_110; 
  assign _T_112 = {_T_111, 2'h0}; 
  assign _T_113 = _T_112[7:0]; 
  assign _T_114 = _T_111 | _T_113; 
  assign _T_115 = {_T_114, 4'h0}; 
  assign _T_116 = _T_115[7:0]; 
  assign _T_117 = _T_114 | _T_116; 
  assign _T_119 = ~ _T_117; 
  assign _GEN_30 = {{1'd0}, _T_107}; 
  assign _T_120 = _GEN_30 | _T_119; 
  assign _T_121 = {_T_94, 1'h0}; 
  assign _T_122 = _T_121[7:0]; 
  assign _T_123 = _T_94 | _T_122; 
  assign _T_124 = {_T_123, 2'h0}; 
  assign _T_125 = _T_124[7:0]; 
  assign _T_126 = _T_123 | _T_125; 
  assign _T_127 = {_T_126, 4'h0}; 
  assign _T_128 = _T_127[7:0]; 
  assign _T_129 = _T_126 | _T_128; 
  assign _T_131 = ~ _T_129; 
  assign _T_132 = _T_120 & _T_131; 
  assign _T_133 = _T_132 & 8'h7; 
  assign _T_86_bits_burst = Queue_1_io_deq_bits_burst; 
  assign _T_134 = _T_86_bits_burst == 2'h0; 
  assign _T_86_bits_size = Queue_1_io_deq_bits_size; 
  assign _T_135 = _T_86_bits_size != 3'h3; 
  assign _T_136 = _T_134 | _T_135; 
  assign _T_137 = _T_136 ? 8'h0 : _T_133; 
  assign _T_138 = {_T_137, 1'h0}; 
  assign _T_139 = _T_138 | 9'h1; 
  assign _T_140 = {1'h0,_T_137}; 
  assign _T_141 = ~ _T_140; 
  assign _T_142 = _T_139 & _T_141; 
  assign _GEN_31 = {{7'd0}, _T_142}; 
  assign _T_143 = _GEN_31 << _T_86_bits_size; 
  assign _GEN_32 = {{16'd0}, _T_143}; 
  assign _T_145 = _T_92 + _GEN_32; 
  assign _T_146 = {_T_86_bits_len,8'hff}; 
  assign _GEN_33 = {{7'd0}, _T_146}; 
  assign _T_147 = _GEN_33 << _T_86_bits_size; 
  assign _T_148 = _T_147[22:8]; 
  assign _T_150 = _T_86_bits_burst == 2'h2; 
  assign _GEN_34 = {{17'd0}, _T_148}; 
  assign _T_151 = _T_145 & _GEN_34; 
  assign _T_152 = ~ _T_86_bits_addr; 
  assign _T_153 = _T_152 | _GEN_34; 
  assign _T_154 = ~ _T_153; 
  assign _T_155 = _T_151 | _T_154; 
  assign _T_157 = _T_137 == _T_91; 
  assign _T_185 = _T_184 == 9'h0; 
  assign _T_179 = _T_185 | _T_172; 
  assign _T_180 = auto_out_awready & _T_179; 
  assign _T_159 = ~ _T_92; 
  assign _T_161 = 10'h7 << _T_86_bits_size; 
  assign _T_162 = _T_161[2:0]; 
  assign _T_163 = ~ _T_162; 
  assign _GEN_36 = {{29'd0}, _T_163}; 
  assign _T_164 = _T_159 | _GEN_36; 
  assign _T_86_valid = Queue_1_io_deq_valid; 
  assign _T_166 = _T_180 & _T_86_valid; 
  assign _T_167 = _T_157 == 1'h0; 
  assign _GEN_37 = {{1'd0}, _T_91}; 
  assign _T_169 = _GEN_37 - _T_142; 
  assign _GEN_9 = _T_166 ? _T_169 : {{1'd0}, _T_90}; 
  assign _T_2_bits_user = Queue_io_deq_bits_user; 
  assign _T_181 = _T_172 == 1'h0; 
  assign _T_182 = _T_86_valid & _T_181; 
  assign _T_175 = _T_182 & _T_185; 
  assign _T_178 = _T_86_valid & _T_179; 
  assign _T_176 = auto_out_awready & _T_178; 
  assign _T_86_bits_user = Queue_1_io_deq_bits_user; 
  assign _T_186 = _T_182 ? _T_142 : 9'h0; 
  assign _T_187 = _T_185 ? _T_186 : _T_184; 
  assign _T_188 = _T_187 == 9'h1; 
  assign _T_170_valid = Queue_2_io_deq_valid; 
  assign _T_199 = _T_185 == 1'h0; 
  assign _T_200 = _T_199 | _T_182; 
  assign _T_201 = _T_170_valid & _T_200; 
  assign _T_189 = auto_out_wready & _T_201; 
  assign _GEN_38 = {{8'd0}, _T_189}; 
  assign _T_191 = _T_187 - _GEN_38; 
  assign _T_193 = _T_189 == 1'h0; 
  assign _T_194 = _T_187 != 9'h0; 
  assign _T_195 = _T_193 | _T_194; 
  assign _T_197 = _T_195 | reset; 
  assign _T_198 = _T_197 == 1'h0; 
  assign _T_205 = _T_201 == 1'h0; 
  assign _T_170_bits_last = Queue_2_io_deq_bits_last; 
  assign _T_206 = _T_170_bits_last == 1'h0; 
  assign _T_207 = _T_205 | _T_206; 
  assign _T_208 = _T_207 | _T_188; 
  assign _T_210 = _T_208 | reset; 
  assign _T_211 = _T_210 == 1'h0; 
  assign _T_212 = auto_out_ruser[0]; 
  assign _T_215 = auto_out_buser[0]; 
  assign _T_217 = _T_215 == 1'h0; 
  assign _T_218 = auto_in_bready | _T_217; 
  assign _GEN_13 = auto_out_bid ? _T_221_1 : _T_221_0; 
  assign _T_224 = 2'h1 << auto_out_bid; 
  assign _T_226 = _T_224[0]; 
  assign _T_227 = _T_224[1]; 
  assign _T_228 = _T_218 & auto_out_bvalid; 
  assign _T_229 = _T_226 & _T_228; 
  assign _T_230 = _T_221_0 | auto_out_bresp; 
  assign _T_233 = _T_227 & _T_228; 
  assign _T_234 = _T_221_1 | auto_out_bresp; 
  assign auto_in_awready = Queue_1_io_enq_ready; 
  assign auto_in_wready = Queue_2_io_enq_ready; 
  assign auto_in_bvalid = auto_out_bvalid & _T_215; 
  assign auto_in_bid = auto_out_bid; 
  assign auto_in_bresp = auto_out_bresp | _GEN_13; 
  assign auto_in_buser = auto_out_buser[16:1]; 
  assign auto_in_arready = Queue_io_enq_ready; 
  assign auto_in_rvalid = auto_out_rvalid; 
  assign auto_in_rid = auto_out_rid; 
  assign auto_in_rdata = auto_out_rdata; 
  assign auto_in_rresp = auto_out_rresp; 
  assign auto_in_ruser = auto_out_ruser[16:1]; 
  assign auto_in_rlast = auto_out_rlast & _T_212; 
  assign auto_out_awvalid = _T_86_valid & _T_179; 
  assign auto_out_awid = Queue_1_io_deq_bits_id; 
  assign auto_out_awaddr = ~ _T_164; 
  assign auto_out_awlen = _T_136 ? 8'h0 : _T_133; 
  assign auto_out_awsize = Queue_1_io_deq_bits_size; 
  assign auto_out_awuser = {_T_86_bits_user,_T_157}; 
  assign auto_out_wvalid = _T_170_valid & _T_200; 
  assign auto_out_wdata = Queue_2_io_deq_bits_data; 
  assign auto_out_wstrb = Queue_2_io_deq_bits_strb; 
  assign auto_out_wlast = _T_187 == 9'h1; 
  assign auto_out_bready = auto_in_bready | _T_217; 
  assign auto_out_arvalid = Queue_io_deq_valid; 
  assign auto_out_arid = Queue_io_deq_bits_id; 
  assign auto_out_araddr = ~ _T_80; 
  assign auto_out_arlen = _T_52 ? 8'h0 : _T_49; 
  assign auto_out_arsize = Queue_io_deq_bits_size; 
  assign auto_out_aruser = {_T_2_bits_user,_T_73}; 
  assign auto_out_rready = auto_in_rready; 
  assign Queue_clock = clock; 
  assign Queue_reset = reset; 
  assign Queue_io_enq_valid = auto_in_arvalid; 
  assign Queue_io_enq_bits_id = auto_in_arid; 
  assign Queue_io_enq_bits_addr = auto_in_araddr; 
  assign Queue_io_enq_bits_len = auto_in_arlen; 
  assign Queue_io_enq_bits_size = auto_in_arsize; 
  assign Queue_io_enq_bits_burst = auto_in_arburst; 
  assign Queue_io_enq_bits_user = auto_in_aruser; 
  assign Queue_io_deq_ready = auto_out_arready & _T_73; 
  assign Queue_1_clock = clock; 
  assign Queue_1_reset = reset; 
  assign Queue_1_io_enq_valid = auto_in_awvalid; 
  assign Queue_1_io_enq_bits_id = auto_in_awid; 
  assign Queue_1_io_enq_bits_addr = auto_in_awaddr; 
  assign Queue_1_io_enq_bits_len = auto_in_awlen; 
  assign Queue_1_io_enq_bits_size = auto_in_awsize; 
  assign Queue_1_io_enq_bits_burst = auto_in_awburst; 
  assign Queue_1_io_enq_bits_user = auto_in_awuser; 
  assign Queue_1_io_deq_ready = _T_180 & _T_157; 
  assign Queue_2_clock = clock; 
  assign Queue_2_reset = reset; 
  assign Queue_2_io_enq_valid = auto_in_wvalid; 
  assign Queue_2_io_enq_bits_data = auto_in_wdata; 
  assign Queue_2_io_enq_bits_strb = auto_in_wstrb; 
  assign Queue_2_io_enq_bits_last = auto_in_wlast; 
  assign Queue_2_io_deq_ready = auto_out_wready & _T_200; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_4 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_5 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_6 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_88 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_89 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_90 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_184 = _RAND_6[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_172 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_221_0 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_221_1 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_4 <= 1'h0;
    end else begin
      if (_T_82) begin
        _T_4 <= _T_83;
      end
    end
    if (_T_82) begin
      if (_T_50) begin
        _T_5 <= _T_2_bits_addr;
      end else begin
        if (_T_66) begin
          _T_5 <= _T_71;
        end else begin
          _T_5 <= _T_61;
        end
      end
    end
    _T_6 <= _GEN_4[7:0];
    if (reset) begin
      _T_88 <= 1'h0;
    end else begin
      if (_T_166) begin
        _T_88 <= _T_167;
      end
    end
    if (_T_166) begin
      if (_T_134) begin
        _T_89 <= _T_86_bits_addr;
      end else begin
        if (_T_150) begin
          _T_89 <= _T_155;
        end else begin
          _T_89 <= _T_145;
        end
      end
    end
    _T_90 <= _GEN_9[7:0];
    if (reset) begin
      _T_184 <= 9'h0;
    end else begin
      _T_184 <= _T_191;
    end
    if (reset) begin
      _T_172 <= 1'h0;
    end else begin
      if (_T_176) begin
        _T_172 <= 1'h0;
      end else begin
        if (_T_175) begin
          _T_172 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_221_0 <= 2'h0;
    end else begin
      if (_T_229) begin
        if (_T_215) begin
          _T_221_0 <= 2'h0;
        end else begin
          _T_221_0 <= _T_230;
        end
      end
    end
    if (reset) begin
      _T_221_1 <= 2'h0;
    end else begin
      if (_T_233) begin
        if (_T_215) begin
          _T_221_1 <= 2'h0;
        end else begin
          _T_221_1 <= _T_234;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_198) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:167 assert (!out.w.fire() || w_todo =/= UInt(0)) // underflow impossible\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_198) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_211) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:176 assert (!out.w.valid || !in_w.bits.last || w_last)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_211) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_AXI4IdIndexer_1( 
  output        auto_in_awready, 
  input         auto_in_awvalid, 
  input  [4:0]  auto_in_awid, 
  input  [30:0] auto_in_awaddr, 
  input  [7:0]  auto_in_awlen, 
  input  [2:0]  auto_in_awsize, 
  input  [1:0]  auto_in_awburst, 
  input         auto_in_awlock, 
  input  [3:0]  auto_in_awcache, 
  input  [2:0]  auto_in_awprot, 
  input  [3:0]  auto_in_awqos, 
  input  [10:0] auto_in_awuser, 
  input  [63:0] auto_in_awinstret, 
  output        auto_in_wready, 
  input         auto_in_wvalid, 
  input  [63:0] auto_in_wdata, 
  input  [7:0]  auto_in_wstrb, 
  input         auto_in_wlast, 
  input         auto_in_bready, 
  output        auto_in_bvalid, 
  output [4:0]  auto_in_bid, 
  output [1:0]  auto_in_bresp, 
  output [10:0] auto_in_buser, 
  output        auto_in_arready, 
  input         auto_in_arvalid, 
  input  [4:0]  auto_in_arid, 
  input  [30:0] auto_in_araddr, 
  input  [7:0]  auto_in_arlen, 
  input  [2:0]  auto_in_arsize, 
  input  [1:0]  auto_in_arburst, 
  input         auto_in_arlock, 
  input  [3:0]  auto_in_arcache, 
  input  [2:0]  auto_in_arprot, 
  input  [3:0]  auto_in_arqos, 
  input  [10:0] auto_in_aruser, 
  input  [63:0] auto_in_arinstret, 
  input         auto_in_rready, 
  output        auto_in_rvalid, 
  output [4:0]  auto_in_rid, 
  output [63:0] auto_in_rdata, 
  output [1:0]  auto_in_rresp, 
  output [10:0] auto_in_ruser, 
  output        auto_in_rlast, 
  input         auto_out_awready, 
  output        auto_out_awvalid, 
  output [30:0] auto_out_awaddr, 
  output [7:0]  auto_out_awlen, 
  output [2:0]  auto_out_awsize, 
  output [1:0]  auto_out_awburst, 
  output        auto_out_awlock, 
  output [3:0]  auto_out_awcache, 
  output [2:0]  auto_out_awprot, 
  output [3:0]  auto_out_awqos, 
  output [15:0] auto_out_awuser, 
  output [63:0] auto_out_awinstret, 
  input         auto_out_wready, 
  output        auto_out_wvalid, 
  output [63:0] auto_out_wdata, 
  output [7:0]  auto_out_wstrb, 
  output        auto_out_wlast, 
  output        auto_out_bready, 
  input         auto_out_bvalid, 
  input  [1:0]  auto_out_bresp, 
  input  [15:0] auto_out_buser, 
  input         auto_out_arready, 
  output        auto_out_arvalid, 
  output [30:0] auto_out_araddr, 
  output [7:0]  auto_out_arlen, 
  output [2:0]  auto_out_arsize, 
  output [1:0]  auto_out_arburst, 
  output        auto_out_arlock, 
  output [3:0]  auto_out_arcache, 
  output [2:0]  auto_out_arprot, 
  output [3:0]  auto_out_arqos, 
  output [15:0] auto_out_aruser, 
  output [63:0] auto_out_arinstret, 
  output        auto_out_rready, 
  input         auto_out_rvalid, 
  input  [63:0] auto_out_rdata, 
  input  [1:0]  auto_out_rresp, 
  input  [15:0] auto_out_ruser, 
  input         auto_out_rlast 
);
  assign auto_in_awready = auto_out_awready; 
  assign auto_in_wready = auto_out_wready; 
  assign auto_in_bvalid = auto_out_bvalid; 
  assign auto_in_bid = auto_out_buser[4:0]; 
  assign auto_in_bresp = auto_out_bresp; 
  assign auto_in_buser = auto_out_buser[15:5]; 
  assign auto_in_arready = auto_out_arready; 
  assign auto_in_rvalid = auto_out_rvalid; 
  assign auto_in_rid = auto_out_ruser[4:0]; 
  assign auto_in_rdata = auto_out_rdata; 
  assign auto_in_rresp = auto_out_rresp; 
  assign auto_in_ruser = auto_out_ruser[15:5]; 
  assign auto_in_rlast = auto_out_rlast; 
  assign auto_out_awvalid = auto_in_awvalid; 
  assign auto_out_awaddr = auto_in_awaddr; 
  assign auto_out_awlen = auto_in_awlen; 
  assign auto_out_awsize = auto_in_awsize; 
  assign auto_out_awburst = auto_in_awburst; 
  assign auto_out_awlock = auto_in_awlock; 
  assign auto_out_awcache = auto_in_awcache; 
  assign auto_out_awprot = auto_in_awprot; 
  assign auto_out_awqos = auto_in_awqos; 
  assign auto_out_awuser = {auto_in_awuser,auto_in_awid}; 
  assign auto_out_awinstret = auto_in_awinstret; 
  assign auto_out_wvalid = auto_in_wvalid; 
  assign auto_out_wdata = auto_in_wdata; 
  assign auto_out_wstrb = auto_in_wstrb; 
  assign auto_out_wlast = auto_in_wlast; 
  assign auto_out_bready = auto_in_bready; 
  assign auto_out_arvalid = auto_in_arvalid; 
  assign auto_out_araddr = auto_in_araddr; 
  assign auto_out_arlen = auto_in_arlen; 
  assign auto_out_arsize = auto_in_arsize; 
  assign auto_out_arburst = auto_in_arburst; 
  assign auto_out_arlock = auto_in_arlock; 
  assign auto_out_arcache = auto_in_arcache; 
  assign auto_out_arprot = auto_in_arprot; 
  assign auto_out_arqos = auto_in_arqos; 
  assign auto_out_aruser = {auto_in_aruser,auto_in_arid}; 
  assign auto_out_arinstret = auto_in_arinstret; 
  assign auto_out_rready = auto_in_rready; 
endmodule
module dual_AXI4IdIndexer_2( 
  output        auto_in_awready, 
  input         auto_in_awvalid, 
  input  [16:0] auto_in_awid, 
  input  [31:0] auto_in_awaddr, 
  input  [7:0]  auto_in_awlen, 
  input  [2:0]  auto_in_awsize, 
  input  [1:0]  auto_in_awburst, 
  output        auto_in_wready, 
  input         auto_in_wvalid, 
  input  [63:0] auto_in_wdata, 
  input  [7:0]  auto_in_wstrb, 
  input         auto_in_wlast, 
  input         auto_in_bready, 
  output        auto_in_bvalid, 
  output [16:0] auto_in_bid, 
  output [1:0]  auto_in_bresp, 
  output        auto_in_arready, 
  input         auto_in_arvalid, 
  input  [16:0] auto_in_arid, 
  input  [31:0] auto_in_araddr, 
  input  [7:0]  auto_in_arlen, 
  input  [2:0]  auto_in_arsize, 
  input  [1:0]  auto_in_arburst, 
  input         auto_in_rready, 
  output        auto_in_rvalid, 
  output [16:0] auto_in_rid, 
  output [63:0] auto_in_rdata, 
  output [1:0]  auto_in_rresp, 
  output        auto_in_rlast, 
  input         auto_out_awready, 
  output        auto_out_awvalid, 
  output        auto_out_awid, 
  output [31:0] auto_out_awaddr, 
  output [7:0]  auto_out_awlen, 
  output [2:0]  auto_out_awsize, 
  output [1:0]  auto_out_awburst, 
  output [15:0] auto_out_awuser, 
  input         auto_out_wready, 
  output        auto_out_wvalid, 
  output [63:0] auto_out_wdata, 
  output [7:0]  auto_out_wstrb, 
  output        auto_out_wlast, 
  output        auto_out_bready, 
  input         auto_out_bvalid, 
  input         auto_out_bid, 
  input  [1:0]  auto_out_bresp, 
  input  [15:0] auto_out_buser, 
  input         auto_out_arready, 
  output        auto_out_arvalid, 
  output        auto_out_arid, 
  output [31:0] auto_out_araddr, 
  output [7:0]  auto_out_arlen, 
  output [2:0]  auto_out_arsize, 
  output [1:0]  auto_out_arburst, 
  output [15:0] auto_out_aruser, 
  output        auto_out_rready, 
  input         auto_out_rvalid, 
  input         auto_out_rid, 
  input  [63:0] auto_out_rdata, 
  input  [1:0]  auto_out_rresp, 
  input  [15:0] auto_out_ruser, 
  input         auto_out_rlast 
);
  assign auto_in_awready = auto_out_awready; 
  assign auto_in_wready = auto_out_wready; 
  assign auto_in_bvalid = auto_out_bvalid; 
  assign auto_in_bid = {auto_out_buser,auto_out_bid}; 
  assign auto_in_bresp = auto_out_bresp; 
  assign auto_in_arready = auto_out_arready; 
  assign auto_in_rvalid = auto_out_rvalid; 
  assign auto_in_rid = {auto_out_ruser,auto_out_rid}; 
  assign auto_in_rdata = auto_out_rdata; 
  assign auto_in_rresp = auto_out_rresp; 
  assign auto_in_rlast = auto_out_rlast; 
  assign auto_out_awvalid = auto_in_awvalid; 
  assign auto_out_awid = auto_in_awid[0]; 
  assign auto_out_awaddr = auto_in_awaddr; 
  assign auto_out_awlen = auto_in_awlen; 
  assign auto_out_awsize = auto_in_awsize; 
  assign auto_out_awburst = auto_in_awburst; 
  assign auto_out_awuser = auto_in_awid[16:1]; 
  assign auto_out_wvalid = auto_in_wvalid; 
  assign auto_out_wdata = auto_in_wdata; 
  assign auto_out_wstrb = auto_in_wstrb; 
  assign auto_out_wlast = auto_in_wlast; 
  assign auto_out_bready = auto_in_bready; 
  assign auto_out_arvalid = auto_in_arvalid; 
  assign auto_out_arid = auto_in_arid[0]; 
  assign auto_out_araddr = auto_in_araddr; 
  assign auto_out_arlen = auto_in_arlen; 
  assign auto_out_arsize = auto_in_arsize; 
  assign auto_out_arburst = auto_in_arburst; 
  assign auto_out_aruser = auto_in_arid[16:1]; 
  assign auto_out_rready = auto_in_rready; 
endmodule
module dual_AXI4IdIndexer( 
  output        auto_in_awready, 
  input         auto_in_awvalid, 
  input  [4:0]  auto_in_awid, 
  input  [31:0] auto_in_awaddr, 
  input  [7:0]  auto_in_awlen, 
  input  [2:0]  auto_in_awsize, 
  input  [1:0]  auto_in_awburst, 
  input         auto_in_awlock, 
  input  [3:0]  auto_in_awcache, 
  input  [2:0]  auto_in_awprot, 
  input  [3:0]  auto_in_awqos, 
  input  [10:0] auto_in_awuser, 
  input  [63:0] auto_in_awinstret, 
  output        auto_in_wready, 
  input         auto_in_wvalid, 
  input  [63:0] auto_in_wdata, 
  input  [7:0]  auto_in_wstrb, 
  input         auto_in_wlast, 
  input         auto_in_bready, 
  output        auto_in_bvalid, 
  output [4:0]  auto_in_bid, 
  output [1:0]  auto_in_bresp, 
  output [10:0] auto_in_buser, 
  output        auto_in_arready, 
  input         auto_in_arvalid, 
  input  [4:0]  auto_in_arid, 
  input  [31:0] auto_in_araddr, 
  input  [7:0]  auto_in_arlen, 
  input  [2:0]  auto_in_arsize, 
  input  [1:0]  auto_in_arburst, 
  input         auto_in_arlock, 
  input  [3:0]  auto_in_arcache, 
  input  [2:0]  auto_in_arprot, 
  input  [3:0]  auto_in_arqos, 
  input  [10:0] auto_in_aruser, 
  input  [63:0] auto_in_arinstret, 
  input         auto_in_rready, 
  output        auto_in_rvalid, 
  output [4:0]  auto_in_rid, 
  output [63:0] auto_in_rdata, 
  output [1:0]  auto_in_rresp, 
  output [10:0] auto_in_ruser, 
  output        auto_in_rlast, 
  input         auto_out_awready, 
  output        auto_out_awvalid, 
  output [3:0]  auto_out_awid, 
  output [31:0] auto_out_awaddr, 
  output [7:0]  auto_out_awlen, 
  output [2:0]  auto_out_awsize, 
  output [1:0]  auto_out_awburst, 
  output        auto_out_awlock, 
  output [3:0]  auto_out_awcache, 
  output [2:0]  auto_out_awprot, 
  output [3:0]  auto_out_awqos, 
  output [11:0] auto_out_awuser, 
  output [63:0] auto_out_awinstret, 
  input         auto_out_wready, 
  output        auto_out_wvalid, 
  output [63:0] auto_out_wdata, 
  output [7:0]  auto_out_wstrb, 
  output        auto_out_wlast, 
  output        auto_out_bready, 
  input         auto_out_bvalid, 
  input  [3:0]  auto_out_bid, 
  input  [1:0]  auto_out_bresp, 
  input  [11:0] auto_out_buser, 
  input         auto_out_arready, 
  output        auto_out_arvalid, 
  output [3:0]  auto_out_arid, 
  output [31:0] auto_out_araddr, 
  output [7:0]  auto_out_arlen, 
  output [2:0]  auto_out_arsize, 
  output [1:0]  auto_out_arburst, 
  output        auto_out_arlock, 
  output [3:0]  auto_out_arcache, 
  output [2:0]  auto_out_arprot, 
  output [3:0]  auto_out_arqos, 
  output [11:0] auto_out_aruser, 
  output [63:0] auto_out_arinstret, 
  output        auto_out_rready, 
  input         auto_out_rvalid, 
  input  [3:0]  auto_out_rid, 
  input  [63:0] auto_out_rdata, 
  input  [1:0]  auto_out_rresp, 
  input  [11:0] auto_out_ruser, 
  input         auto_out_rlast 
);
  wire  _T_2; 
  wire  _T_4; 
  wire [15:0] _T_8; 
  wire [15:0] _T_9; 
  assign _T_2 = auto_in_arid[4:4]; 
  assign _T_4 = auto_in_awid[4:4]; 
  assign _T_8 = {auto_out_ruser,auto_out_rid}; 
  assign _T_9 = {auto_out_buser,auto_out_bid}; 
  assign auto_in_awready = auto_out_awready; 
  assign auto_in_wready = auto_out_wready; 
  assign auto_in_bvalid = auto_out_bvalid; 
  assign auto_in_bid = _T_9[4:0]; 
  assign auto_in_bresp = auto_out_bresp; 
  assign auto_in_buser = auto_out_buser[11:1]; 
  assign auto_in_arready = auto_out_arready; 
  assign auto_in_rvalid = auto_out_rvalid; 
  assign auto_in_rid = _T_8[4:0]; 
  assign auto_in_rdata = auto_out_rdata; 
  assign auto_in_rresp = auto_out_rresp; 
  assign auto_in_ruser = auto_out_ruser[11:1]; 
  assign auto_in_rlast = auto_out_rlast; 
  assign auto_out_awvalid = auto_in_awvalid; 
  assign auto_out_awid = auto_in_awid[3:0]; 
  assign auto_out_awaddr = auto_in_awaddr; 
  assign auto_out_awlen = auto_in_awlen; 
  assign auto_out_awsize = auto_in_awsize; 
  assign auto_out_awburst = auto_in_awburst; 
  assign auto_out_awlock = auto_in_awlock; 
  assign auto_out_awcache = auto_in_awcache; 
  assign auto_out_awprot = auto_in_awprot; 
  assign auto_out_awqos = auto_in_awqos; 
  assign auto_out_awuser = {auto_in_awuser,_T_4}; 
  assign auto_out_awinstret = auto_in_awinstret; 
  assign auto_out_wvalid = auto_in_wvalid; 
  assign auto_out_wdata = auto_in_wdata; 
  assign auto_out_wstrb = auto_in_wstrb; 
  assign auto_out_wlast = auto_in_wlast; 
  assign auto_out_bready = auto_in_bready; 
  assign auto_out_arvalid = auto_in_arvalid; 
  assign auto_out_arid = auto_in_arid[3:0]; 
  assign auto_out_araddr = auto_in_araddr; 
  assign auto_out_arlen = auto_in_arlen; 
  assign auto_out_arsize = auto_in_arsize; 
  assign auto_out_arburst = auto_in_arburst; 
  assign auto_out_arlock = auto_in_arlock; 
  assign auto_out_arcache = auto_in_arcache; 
  assign auto_out_arprot = auto_in_arprot; 
  assign auto_out_arqos = auto_in_arqos; 
  assign auto_out_aruser = {auto_in_aruser,_T_2}; 
  assign auto_out_arinstret = auto_in_arinstret; 
  assign auto_out_rready = auto_in_rready; 
endmodule
module dual_AXI4ToTL_top( 
  input         clock, 
  input         reset, 
  output        auto_in_awready, 
  input         auto_in_awvalid, 
  input         auto_in_awid, 
  input  [31:0] auto_in_awaddr, 
  input  [7:0]  auto_in_awlen, 
  input  [2:0]  auto_in_awsize, 
  output        auto_in_wready, 
  input         auto_in_wvalid, 
  input  [63:0] auto_in_wdata, 
  input  [7:0]  auto_in_wstrb, 
  input         auto_in_wlast, 
  input         auto_in_bready, 
  output        auto_in_bvalid, 
  output        auto_in_bid, 
  output [1:0]  auto_in_bresp, 
  output        auto_in_arready, 
  input         auto_in_arvalid, 
  input         auto_in_arid, 
  input  [31:0] auto_in_araddr, 
  input  [7:0]  auto_in_arlen, 
  input  [2:0]  auto_in_arsize, 
  input         auto_in_rready, 
  output        auto_in_rvalid, 
  output        auto_in_rid, 
  output [63:0] auto_in_rdata, 
  output [1:0]  auto_in_rresp, 
  output        auto_in_rlast, 
  input         auto_out_a_ready, 
  output        auto_out_a_valid, 
  output [2:0]  auto_out_a_bits_opcode, 
  output [2:0]  auto_out_a_bits_param, 
  output [2:0]  auto_out_a_bits_size, 
  output [2:0]  auto_out_a_bits_source, 
  output [31:0] auto_out_a_bits_address, 
  output [7:0]  auto_out_a_bits_mask, 
  output [63:0] auto_out_a_bits_data, 
  output        auto_out_a_bits_corrupt, 
  output        auto_out_d_ready, 
  input         auto_out_d_valid, 
  input  [2:0]  auto_out_d_bits_opcode, 
  input  [2:0]  auto_out_d_bits_size, 
  input  [2:0]  auto_out_d_bits_source, 
  input         auto_out_d_bits_denied, 
  input  [63:0] auto_out_d_bits_data, 
  input         auto_out_d_bits_corrupt 
);
  wire  Queue_clock; 
  wire  Queue_reset; 
  wire  Queue_io_enq_ready; 
  wire  Queue_io_enq_valid; 
  wire  Queue_io_enq_bits_id; 
  wire [63:0] Queue_io_enq_bits_data; 
  wire [1:0] Queue_io_enq_bits_resp; 
  wire  Queue_io_enq_bits_last; 
  wire  Queue_io_deq_ready; 
  wire  Queue_io_deq_valid; 
  wire  Queue_io_deq_bits_id; 
  wire [63:0] Queue_io_deq_bits_data; 
  wire [1:0] Queue_io_deq_bits_resp; 
  wire  Queue_io_deq_bits_last; 
  wire  Queue_1_clock; 
  wire  Queue_1_reset; 
  wire  Queue_1_io_enq_ready; 
  wire  Queue_1_io_enq_valid; 
  wire  Queue_1_io_enq_bits_id; 
  wire [1:0] Queue_1_io_enq_bits_resp; 
  wire  Queue_1_io_deq_ready; 
  wire  Queue_1_io_deq_valid; 
  wire  Queue_1_io_deq_bits_id; 
  wire [1:0] Queue_1_io_deq_bits_resp; 
  wire [15:0] _T_3; 
  wire [22:0] _GEN_16; 
  wire [22:0] _T_4; 
  wire [14:0] _T_5; 
  wire [15:0] _T_6; 
  wire [15:0] _T_7; 
  wire [15:0] _T_8; 
  wire [15:0] _T_9; 
  wire [15:0] _T_10; 
  wire [7:0] _T_11; 
  wire [7:0] _T_12; 
  wire  _T_13; 
  wire [7:0] _T_14; 
  wire [3:0] _T_15; 
  wire [3:0] _T_16; 
  wire  _T_17; 
  wire [3:0] _T_18; 
  wire [1:0] _T_19; 
  wire [1:0] _T_20; 
  wire  _T_21; 
  wire [1:0] _T_22; 
  wire  _T_23; 
  wire [3:0] _T_26; 
  wire  _T_28; 
  wire [31:0] _T_31; 
  wire [32:0] _T_32; 
  wire [32:0] _T_33; 
  wire [32:0] _T_34; 
  wire  _T_35; 
  wire [31:0] _T_36; 
  wire [32:0] _T_37; 
  wire [32:0] _T_38; 
  wire [32:0] _T_39; 
  wire  _T_40; 
  wire [31:0] _T_41; 
  wire [32:0] _T_42; 
  wire [32:0] _T_43; 
  wire [32:0] _T_44; 
  wire  _T_45; 
  wire  _T_46; 
  wire  _T_47; 
  wire  _T_48; 
  wire [2:0] _T_50; 
  wire [28:0] _GEN_17; 
  wire [28:0] _T_51; 
  wire [31:0] _T_52; 
  reg [1:0] _T_54_0; 
  reg [31:0] _RAND_0;
  reg [1:0] _T_54_1; 
  reg [31:0] _RAND_1;
  wire [1:0] _GEN_1; 
  wire  _T_55; 
  wire  _T_58; 
  wire [29:0] _T_60; 
  wire [14:0] _T_61; 
  wire [14:0] _T_62; 
  wire  _T_63; 
  wire  _T_64; 
  wire  _T_66; 
  wire  _T_67; 
  wire [1:0] _T_81; 
  wire [3:0] _T_82; 
  wire [2:0] _T_83; 
  wire [2:0] _T_84; 
  wire  _T_85; 
  wire  _T_86; 
  wire  _T_87; 
  wire  _T_88; 
  wire  _T_90; 
  wire  _T_91; 
  wire  _T_93; 
  wire  _T_94; 
  wire  _T_95; 
  wire  _T_96; 
  wire  _T_97; 
  wire  _T_98; 
  wire  _T_99; 
  wire  _T_100; 
  wire  _T_101; 
  wire  _T_102; 
  wire  _T_103; 
  wire  _T_104; 
  wire  _T_105; 
  wire  _T_106; 
  wire  _T_107; 
  wire  _T_108; 
  wire  _T_109; 
  wire  _T_110; 
  wire  _T_111; 
  wire  _T_112; 
  wire  _T_113; 
  wire  _T_114; 
  wire  _T_115; 
  wire  _T_116; 
  wire  _T_117; 
  wire  _T_118; 
  wire  _T_119; 
  wire  _T_120; 
  wire  _T_121; 
  wire  _T_122; 
  wire  _T_123; 
  wire  _T_124; 
  wire  _T_125; 
  wire  _T_126; 
  wire  _T_127; 
  wire  _T_128; 
  wire  _T_129; 
  wire  _T_130; 
  wire  _T_131; 
  wire  _T_132; 
  wire  _T_133; 
  wire  _T_134; 
  wire  _T_135; 
  wire  _T_136; 
  wire [1:0] _T_145; 
  wire  _T_147; 
  wire  _T_148; 
  reg [7:0] _T_260; 
  reg [31:0] _RAND_2;
  wire  _T_261; 
  wire  _T_234; 
  wire [1:0] _T_263; 
  reg [1:0] _T_270; 
  reg [31:0] _RAND_3;
  wire [1:0] _T_271; 
  wire [1:0] _T_272; 
  wire [3:0] _T_273; 
  wire [2:0] _T_274; 
  wire [3:0] _GEN_18; 
  wire [3:0] _T_275; 
  wire [2:0] _T_277; 
  wire [3:0] _T_278; 
  wire [3:0] _GEN_19; 
  wire [3:0] _T_279; 
  wire [1:0] _T_280; 
  wire [1:0] _T_281; 
  wire [1:0] _T_282; 
  wire [1:0] _T_283; 
  wire  _T_292; 
  reg  _T_325_0; 
  reg [31:0] _RAND_4;
  wire  _T_327_0; 
  wire  _T_328; 
  wire  _T_149; 
  wire  _T_150; 
  wire [1:0] _T_152; 
  wire  _T_154; 
  wire [1:0] _T_156; 
  wire [15:0] _T_158; 
  wire [22:0] _GEN_20; 
  wire [22:0] _T_159; 
  wire [14:0] _T_160; 
  wire [15:0] _T_161; 
  wire [15:0] _T_162; 
  wire [15:0] _T_163; 
  wire [15:0] _T_164; 
  wire [15:0] _T_165; 
  wire [7:0] _T_166; 
  wire [7:0] _T_167; 
  wire  _T_168; 
  wire [7:0] _T_169; 
  wire [3:0] _T_170; 
  wire [3:0] _T_171; 
  wire  _T_172; 
  wire [3:0] _T_173; 
  wire [1:0] _T_174; 
  wire [1:0] _T_175; 
  wire  _T_176; 
  wire [1:0] _T_177; 
  wire  _T_178; 
  wire [3:0] _T_181; 
  wire  _T_183; 
  wire [31:0] _T_186; 
  wire [32:0] _T_187; 
  wire [32:0] _T_188; 
  wire [32:0] _T_189; 
  wire  _T_190; 
  wire [31:0] _T_191; 
  wire [32:0] _T_192; 
  wire [32:0] _T_193; 
  wire [32:0] _T_194; 
  wire  _T_195; 
  wire [31:0] _T_196; 
  wire [32:0] _T_197; 
  wire [32:0] _T_198; 
  wire [32:0] _T_199; 
  wire  _T_200; 
  wire  _T_201; 
  wire  _T_202; 
  wire  _T_203; 
  wire [2:0] _T_205; 
  wire [28:0] _GEN_21; 
  wire [28:0] _T_206; 
  wire [31:0] _T_207; 
  reg [1:0] _T_209_0; 
  reg [31:0] _RAND_5;
  reg [1:0] _T_209_1; 
  reg [31:0] _RAND_6;
  wire [1:0] _GEN_5; 
  wire  _T_210; 
  wire  _T_213; 
  wire [29:0] _T_215; 
  wire [14:0] _T_216; 
  wire [14:0] _T_217; 
  wire  _T_218; 
  wire  _T_219; 
  wire  _T_221; 
  wire  _T_222; 
  wire  _T_224; 
  wire  _T_225; 
  wire  _T_226; 
  wire  _T_227; 
  wire  _T_229; 
  wire  _T_230; 
  wire  _T_293; 
  reg  _T_325_1; 
  reg [31:0] _RAND_7;
  wire  _T_327_1; 
  wire  _T_329; 
  wire  _T_231; 
  wire  _T_232; 
  wire [1:0] _T_248; 
  wire  _T_250; 
  wire  _T_251; 
  wire  _T_252; 
  wire  _T_253; 
  wire [1:0] _T_255; 
  wire  _T_257; 
  wire [1:0] _T_259; 
  wire  _T_262; 
  wire  _T_265; 
  wire  _T_267; 
  wire  _T_268; 
  wire  _T_284; 
  wire  _T_285; 
  wire [1:0] _T_286; 
  wire [2:0] _T_287; 
  wire [1:0] _T_288; 
  wire [1:0] _T_289; 
  wire  _T_295; 
  wire  _T_296; 
  wire  _T_299; 
  wire  _T_301; 
  wire  _T_304; 
  wire  _T_305; 
  wire  _T_308; 
  wire  _T_309; 
  wire  _T_310; 
  wire  _T_311; 
  wire  _T_313; 
  wire  _T_315; 
  wire  _T_316; 
  wire  _T_331; 
  wire  _T_332; 
  wire  _T_333; 
  wire  _T_335; 
  wire  _T_320; 
  wire [7:0] _GEN_22; 
  wire [7:0] _T_322; 
  wire  _T_326_0; 
  wire  _T_326_1; 
  wire [141:0] _T_339; 
  wire [2:0] _T_79_size; 
  wire [185:0] _T_344; 
  wire [185:0] _T_345; 
  wire [2:0] _T_246_size; 
  wire [185:0] _T_354; 
  wire [185:0] _T_355; 
  wire [185:0] _T_356; 
  wire  _T_371; 
  wire  _T_373; 
  wire  _T_370_ready; 
  wire  _T_369_ready; 
  wire  _T_393; 
  wire  _T_374; 
  wire [12:0] _T_376; 
  wire [5:0] _T_377; 
  wire [5:0] _T_378; 
  wire [2:0] _T_379; 
  wire [2:0] _T_381; 
  reg [2:0] _T_382; 
  reg [31:0] _RAND_8;
  wire [2:0] _T_384; 
  wire  _T_385; 
  wire  _T_386; 
  wire  _T_387; 
  wire  _T_395; 
  reg [1:0] _T_402_0; 
  reg [31:0] _RAND_9;
  reg [1:0] _T_402_1; 
  reg [31:0] _RAND_10;
  wire  _T_400_bits_id; 
  wire [1:0] _GEN_11; 
  wire [1:0] _GEN_13; 
  wire  _T_403; 
  wire [1:0] _T_405; 
  wire  _T_407; 
  wire  _T_408; 
  wire  _T_400_valid; 
  wire  _T_417; 
  wire  _T_409; 
  wire  _T_410; 
  wire [1:0] _T_412; 
  wire  _T_414; 
  wire [1:0] _T_416; 
  dual_Queue_58 dual_Queue ( 
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_resp(Queue_io_enq_bits_resp),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_resp(Queue_io_deq_bits_resp),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  dual_Queue_59 Queue_1 ( 
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_id(Queue_1_io_enq_bits_id),
    .io_enq_bits_resp(Queue_1_io_enq_bits_resp),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_id(Queue_1_io_deq_bits_id),
    .io_deq_bits_resp(Queue_1_io_deq_bits_resp)
  );
  assign _T_3 = {auto_in_arlen,8'hff}; 
  assign _GEN_16 = {{7'd0}, _T_3}; 
  assign _T_4 = _GEN_16 << auto_in_arsize; 
  assign _T_5 = _T_4[22:8]; 
  assign _T_6 = {_T_5, 1'h0}; 
  assign _T_7 = _T_6 | 16'h1; 
  assign _T_8 = {1'h0,_T_5}; 
  assign _T_9 = ~ _T_8; 
  assign _T_10 = _T_7 & _T_9; 
  assign _T_11 = _T_10[15:8]; 
  assign _T_12 = _T_10[7:0]; 
  assign _T_13 = _T_11 != 8'h0; 
  assign _T_14 = _T_11 | _T_12; 
  assign _T_15 = _T_14[7:4]; 
  assign _T_16 = _T_14[3:0]; 
  assign _T_17 = _T_15 != 4'h0; 
  assign _T_18 = _T_15 | _T_16; 
  assign _T_19 = _T_18[3:2]; 
  assign _T_20 = _T_18[1:0]; 
  assign _T_21 = _T_19 != 2'h0; 
  assign _T_22 = _T_19 | _T_20; 
  assign _T_23 = _T_22[1]; 
  assign _T_26 = {_T_13,_T_17,_T_21,_T_23}; 
  assign _T_28 = _T_26 <= 4'h6; 
  assign _T_31 = auto_in_araddr ^ 32'h40000000; 
  assign _T_32 = {1'b0,$signed(_T_31)}; 
  assign _T_33 = $signed(_T_32) & $signed(-33'sh20000000); 
  assign _T_34 = $signed(_T_33); 
  assign _T_35 = $signed(_T_34) == $signed(33'sh0); 
  assign _T_36 = auto_in_araddr ^ 32'h80000000; 
  assign _T_37 = {1'b0,$signed(_T_36)}; 
  assign _T_38 = $signed(_T_37) & $signed(-33'sh80000000); 
  assign _T_39 = $signed(_T_38); 
  assign _T_40 = $signed(_T_39) == $signed(33'sh0); 
  assign _T_41 = auto_in_araddr ^ 32'h10000000; 
  assign _T_42 = {1'b0,$signed(_T_41)}; 
  assign _T_43 = $signed(_T_42) & $signed(-33'sh10000000); 
  assign _T_44 = $signed(_T_43); 
  assign _T_45 = $signed(_T_44) == $signed(33'sh0); 
  assign _T_46 = _T_35 | _T_40; 
  assign _T_47 = _T_46 | _T_45; 
  assign _T_48 = _T_28 & _T_47; 
  assign _T_50 = auto_in_araddr[2:0]; 
  assign _GEN_17 = {{26'd0}, _T_50}; 
  assign _T_51 = 29'h10000000 | _GEN_17; 
  assign _T_52 = _T_48 ? auto_in_araddr : {{3'd0}, _T_51}; 
  assign _GEN_1 = auto_in_arid ? _T_54_1 : _T_54_0; 
  assign _T_55 = _GEN_1[0]; 
  assign _T_58 = auto_in_arvalid == 1'h0; 
  assign _T_60 = 30'h7fff << _T_26; 
  assign _T_61 = _T_60[14:0]; 
  assign _T_62 = ~ _T_61; 
  assign _T_63 = _T_5 == _T_62; 
  assign _T_64 = _T_58 | _T_63; 
  assign _T_66 = _T_64 | reset; 
  assign _T_67 = _T_66 == 1'h0; 
  assign _T_81 = _T_26[1:0]; 
  assign _T_82 = 4'h1 << _T_81; 
  assign _T_83 = _T_82[2:0]; 
  assign _T_84 = _T_83 | 3'h1; 
  assign _T_85 = _T_26 >= 4'h3; 
  assign _T_86 = _T_84[2]; 
  assign _T_87 = _T_52[2]; 
  assign _T_88 = _T_87 == 1'h0; 
  assign _T_90 = _T_86 & _T_88; 
  assign _T_91 = _T_85 | _T_90; 
  assign _T_93 = _T_86 & _T_87; 
  assign _T_94 = _T_85 | _T_93; 
  assign _T_95 = _T_84[1]; 
  assign _T_96 = _T_52[1]; 
  assign _T_97 = _T_96 == 1'h0; 
  assign _T_98 = _T_88 & _T_97; 
  assign _T_99 = _T_95 & _T_98; 
  assign _T_100 = _T_91 | _T_99; 
  assign _T_101 = _T_88 & _T_96; 
  assign _T_102 = _T_95 & _T_101; 
  assign _T_103 = _T_91 | _T_102; 
  assign _T_104 = _T_87 & _T_97; 
  assign _T_105 = _T_95 & _T_104; 
  assign _T_106 = _T_94 | _T_105; 
  assign _T_107 = _T_87 & _T_96; 
  assign _T_108 = _T_95 & _T_107; 
  assign _T_109 = _T_94 | _T_108; 
  assign _T_110 = _T_84[0]; 
  assign _T_111 = _T_52[0]; 
  assign _T_112 = _T_111 == 1'h0; 
  assign _T_113 = _T_98 & _T_112; 
  assign _T_114 = _T_110 & _T_113; 
  assign _T_115 = _T_100 | _T_114; 
  assign _T_116 = _T_98 & _T_111; 
  assign _T_117 = _T_110 & _T_116; 
  assign _T_118 = _T_100 | _T_117; 
  assign _T_119 = _T_101 & _T_112; 
  assign _T_120 = _T_110 & _T_119; 
  assign _T_121 = _T_103 | _T_120; 
  assign _T_122 = _T_101 & _T_111; 
  assign _T_123 = _T_110 & _T_122; 
  assign _T_124 = _T_103 | _T_123; 
  assign _T_125 = _T_104 & _T_112; 
  assign _T_126 = _T_110 & _T_125; 
  assign _T_127 = _T_106 | _T_126; 
  assign _T_128 = _T_104 & _T_111; 
  assign _T_129 = _T_110 & _T_128; 
  assign _T_130 = _T_106 | _T_129; 
  assign _T_131 = _T_107 & _T_112; 
  assign _T_132 = _T_110 & _T_131; 
  assign _T_133 = _T_109 | _T_132; 
  assign _T_134 = _T_107 & _T_111; 
  assign _T_135 = _T_110 & _T_134; 
  assign _T_136 = _T_109 | _T_135; 
  assign _T_145 = 2'h1 << auto_in_arid; 
  assign _T_147 = _T_145[0]; 
  assign _T_148 = _T_145[1]; 
  assign _T_261 = _T_260 == 8'h0; 
  assign _T_234 = auto_in_awvalid & auto_in_wvalid; 
  assign _T_263 = {_T_234,auto_in_arvalid}; 
  assign _T_271 = ~ _T_270; 
  assign _T_272 = _T_263 & _T_271; 
  assign _T_273 = {_T_272,_T_234,auto_in_arvalid}; 
  assign _T_274 = _T_273[3:1]; 
  assign _GEN_18 = {{1'd0}, _T_274}; 
  assign _T_275 = _T_273 | _GEN_18; 
  assign _T_277 = _T_275[3:1]; 
  assign _T_278 = {_T_270, 2'h0}; 
  assign _GEN_19 = {{1'd0}, _T_277}; 
  assign _T_279 = _GEN_19 | _T_278; 
  assign _T_280 = _T_279[3:2]; 
  assign _T_281 = _T_279[1:0]; 
  assign _T_282 = _T_280 & _T_281; 
  assign _T_283 = ~ _T_282; 
  assign _T_292 = _T_283[0]; 
  assign _T_327_0 = _T_261 ? _T_292 : _T_325_0; 
  assign _T_328 = auto_out_a_ready & _T_327_0; 
  assign _T_149 = _T_328 & auto_in_arvalid; 
  assign _T_150 = _T_149 & _T_147; 
  assign _T_152 = _T_54_0 + 2'h1; 
  assign _T_154 = _T_149 & _T_148; 
  assign _T_156 = _T_54_1 + 2'h1; 
  assign _T_158 = {auto_in_awlen,8'hff}; 
  assign _GEN_20 = {{7'd0}, _T_158}; 
  assign _T_159 = _GEN_20 << auto_in_awsize; 
  assign _T_160 = _T_159[22:8]; 
  assign _T_161 = {_T_160, 1'h0}; 
  assign _T_162 = _T_161 | 16'h1; 
  assign _T_163 = {1'h0,_T_160}; 
  assign _T_164 = ~ _T_163; 
  assign _T_165 = _T_162 & _T_164; 
  assign _T_166 = _T_165[15:8]; 
  assign _T_167 = _T_165[7:0]; 
  assign _T_168 = _T_166 != 8'h0; 
  assign _T_169 = _T_166 | _T_167; 
  assign _T_170 = _T_169[7:4]; 
  assign _T_171 = _T_169[3:0]; 
  assign _T_172 = _T_170 != 4'h0; 
  assign _T_173 = _T_170 | _T_171; 
  assign _T_174 = _T_173[3:2]; 
  assign _T_175 = _T_173[1:0]; 
  assign _T_176 = _T_174 != 2'h0; 
  assign _T_177 = _T_174 | _T_175; 
  assign _T_178 = _T_177[1]; 
  assign _T_181 = {_T_168,_T_172,_T_176,_T_178}; 
  assign _T_183 = _T_181 <= 4'h6; 
  assign _T_186 = auto_in_awaddr ^ 32'h40000000; 
  assign _T_187 = {1'b0,$signed(_T_186)}; 
  assign _T_188 = $signed(_T_187) & $signed(-33'sh20000000); 
  assign _T_189 = $signed(_T_188); 
  assign _T_190 = $signed(_T_189) == $signed(33'sh0); 
  assign _T_191 = auto_in_awaddr ^ 32'h80000000; 
  assign _T_192 = {1'b0,$signed(_T_191)}; 
  assign _T_193 = $signed(_T_192) & $signed(-33'sh80000000); 
  assign _T_194 = $signed(_T_193); 
  assign _T_195 = $signed(_T_194) == $signed(33'sh0); 
  assign _T_196 = auto_in_awaddr ^ 32'h10000000; 
  assign _T_197 = {1'b0,$signed(_T_196)}; 
  assign _T_198 = $signed(_T_197) & $signed(-33'sh10000000); 
  assign _T_199 = $signed(_T_198); 
  assign _T_200 = $signed(_T_199) == $signed(33'sh0); 
  assign _T_201 = _T_190 | _T_195; 
  assign _T_202 = _T_201 | _T_200; 
  assign _T_203 = _T_183 & _T_202; 
  assign _T_205 = auto_in_awaddr[2:0]; 
  assign _GEN_21 = {{26'd0}, _T_205}; 
  assign _T_206 = 29'h10000000 | _GEN_21; 
  assign _T_207 = _T_203 ? auto_in_awaddr : {{3'd0}, _T_206}; 
  assign _GEN_5 = auto_in_awid ? _T_209_1 : _T_209_0; 
  assign _T_210 = _GEN_5[0]; 
  assign _T_213 = auto_in_awvalid == 1'h0; 
  assign _T_215 = 30'h7fff << _T_181; 
  assign _T_216 = _T_215[14:0]; 
  assign _T_217 = ~ _T_216; 
  assign _T_218 = _T_160 == _T_217; 
  assign _T_219 = _T_213 | _T_218; 
  assign _T_221 = _T_219 | reset; 
  assign _T_222 = _T_221 == 1'h0; 
  assign _T_224 = auto_in_awlen == 8'h0; 
  assign _T_225 = _T_213 | _T_224; 
  assign _T_226 = auto_in_awsize == 3'h3; 
  assign _T_227 = _T_225 | _T_226; 
  assign _T_229 = _T_227 | reset; 
  assign _T_230 = _T_229 == 1'h0; 
  assign _T_293 = _T_283[1]; 
  assign _T_327_1 = _T_261 ? _T_293 : _T_325_1; 
  assign _T_329 = auto_out_a_ready & _T_327_1; 
  assign _T_231 = _T_329 & auto_in_wvalid; 
  assign _T_232 = _T_231 & auto_in_wlast; 
  assign _T_248 = 2'h1 << auto_in_awid; 
  assign _T_250 = _T_248[0]; 
  assign _T_251 = _T_248[1]; 
  assign _T_252 = _T_232 & auto_in_awvalid; 
  assign _T_253 = _T_252 & _T_250; 
  assign _T_255 = _T_209_0 + 2'h1; 
  assign _T_257 = _T_252 & _T_251; 
  assign _T_259 = _T_209_1 + 2'h1; 
  assign _T_262 = _T_261 & auto_out_a_ready; 
  assign _T_265 = _T_263 == _T_263; 
  assign _T_267 = _T_265 | reset; 
  assign _T_268 = _T_267 == 1'h0; 
  assign _T_284 = _T_263 != 2'h0; 
  assign _T_285 = _T_262 & _T_284; 
  assign _T_286 = _T_283 & _T_263; 
  assign _T_287 = {_T_286, 1'h0}; 
  assign _T_288 = _T_287[1:0]; 
  assign _T_289 = _T_286 | _T_288; 
  assign _T_295 = _T_292 & auto_in_arvalid; 
  assign _T_296 = _T_293 & _T_234; 
  assign _T_299 = _T_295 | _T_296; 
  assign _T_301 = _T_295 == 1'h0; 
  assign _T_304 = _T_296 == 1'h0; 
  assign _T_305 = _T_301 | _T_304; 
  assign _T_308 = _T_305 | reset; 
  assign _T_309 = _T_308 == 1'h0; 
  assign _T_310 = auto_in_arvalid | _T_234; 
  assign _T_311 = _T_310 == 1'h0; 
  assign _T_313 = _T_311 | _T_299; 
  assign _T_315 = _T_313 | reset; 
  assign _T_316 = _T_315 == 1'h0; 
  assign _T_331 = _T_325_0 ? auto_in_arvalid : 1'h0; 
  assign _T_332 = _T_325_1 ? _T_234 : 1'h0; 
  assign _T_333 = _T_331 | _T_332; 
  assign _T_335 = _T_261 ? _T_310 : _T_333; 
  assign _T_320 = auto_out_a_ready & _T_335; 
  assign _GEN_22 = {{7'd0}, _T_320}; 
  assign _T_322 = _T_260 - _GEN_22; 
  assign _T_326_0 = _T_261 ? _T_295 : _T_325_0; 
  assign _T_326_1 = _T_261 ? _T_296 : _T_325_1; 
  assign _T_339 = {69'h0,_T_136,_T_133,_T_130,_T_127,_T_124,_T_121,_T_118,_T_115,65'h0}; 
  assign _T_79_size = _T_26[2:0]; 
  assign _T_344 = {6'h20,_T_79_size,auto_in_arid,_T_55,1'h0,_T_52,_T_339}; 
  assign _T_345 = _T_326_0 ? _T_344 : 186'h0; 
  assign _T_246_size = _T_181[2:0]; 
  assign _T_354 = {6'h8,_T_246_size,auto_in_awid,_T_210,1'h1,_T_207,69'h0,auto_in_wstrb,auto_in_wdata,1'h0}; 
  assign _T_355 = _T_326_1 ? _T_354 : 186'h0; 
  assign _T_356 = _T_345 | _T_355; 
  assign _T_371 = auto_out_d_bits_denied | auto_out_d_bits_corrupt; 
  assign _T_373 = auto_out_d_bits_opcode[0]; 
  assign _T_370_ready = Queue_io_enq_ready; 
  assign _T_369_ready = Queue_1_io_enq_ready; 
  assign _T_393 = _T_373 ? _T_370_ready : _T_369_ready; 
  assign _T_374 = _T_393 & auto_out_d_valid; 
  assign _T_376 = 13'h3f << auto_out_d_bits_size; 
  assign _T_377 = _T_376[5:0]; 
  assign _T_378 = ~ _T_377; 
  assign _T_379 = _T_378[5:3]; 
  assign _T_381 = _T_373 ? _T_379 : 3'h0; 
  assign _T_384 = _T_382 - 3'h1; 
  assign _T_385 = _T_382 == 3'h0; 
  assign _T_386 = _T_382 == 3'h1; 
  assign _T_387 = _T_381 == 3'h0; 
  assign _T_395 = _T_373 == 1'h0; 
  assign _T_400_bits_id = Queue_1_io_deq_bits_id; 
  assign _GEN_11 = _T_400_bits_id ? _T_402_1 : _T_402_0; 
  assign _GEN_13 = _T_400_bits_id ? _T_209_1 : _T_209_0; 
  assign _T_403 = _GEN_11 != _GEN_13; 
  assign _T_405 = 2'h1 << _T_400_bits_id; 
  assign _T_407 = _T_405[0]; 
  assign _T_408 = _T_405[1]; 
  assign _T_400_valid = Queue_1_io_deq_valid; 
  assign _T_417 = _T_400_valid & _T_403; 
  assign _T_409 = auto_in_bready & _T_417; 
  assign _T_410 = _T_409 & _T_407; 
  assign _T_412 = _T_402_0 + 2'h1; 
  assign _T_414 = _T_409 & _T_408; 
  assign _T_416 = _T_402_1 + 2'h1; 
  assign auto_in_awready = _T_231 & auto_in_wlast; 
  assign auto_in_wready = _T_329 & auto_in_awvalid; 
  assign auto_in_bvalid = _T_400_valid & _T_403; 
  assign auto_in_bid = Queue_1_io_deq_bits_id; 
  assign auto_in_bresp = Queue_1_io_deq_bits_resp; 
  assign auto_in_arready = auto_out_a_ready & _T_327_0; 
  assign auto_in_rvalid = Queue_io_deq_valid; 
  assign auto_in_rid = Queue_io_deq_bits_id; 
  assign auto_in_rdata = Queue_io_deq_bits_data; 
  assign auto_in_rresp = Queue_io_deq_bits_resp; 
  assign auto_in_rlast = Queue_io_deq_bits_last; 
  assign auto_out_a_valid = _T_261 ? _T_310 : _T_333; 
  assign auto_out_a_bits_opcode = _T_356[185:183]; 
  assign auto_out_a_bits_param = _T_356[182:180]; 
  assign auto_out_a_bits_size = _T_356[179:177]; 
  assign auto_out_a_bits_source = _T_356[176:174]; 
  assign auto_out_a_bits_address = _T_356[173:142]; 
  assign auto_out_a_bits_mask = _T_356[72:65]; 
  assign auto_out_a_bits_data = _T_356[64:1]; 
  assign auto_out_a_bits_corrupt = _T_356[0]; 
  assign auto_out_d_ready = _T_373 ? _T_370_ready : _T_369_ready; 
  assign Queue_clock = clock; 
  assign Queue_reset = reset; 
  assign Queue_io_enq_valid = auto_out_d_valid & _T_373; 
  assign Queue_io_enq_bits_id = auto_out_d_bits_source[2:2]; 
  assign Queue_io_enq_bits_data = auto_out_d_bits_data; 
  assign Queue_io_enq_bits_resp = _T_371 ? 2'h2 : 2'h0; 
  assign Queue_io_enq_bits_last = _T_386 | _T_387; 
  assign Queue_io_deq_ready = auto_in_rready; 
  assign Queue_1_clock = clock; 
  assign Queue_1_reset = reset; 
  assign Queue_1_io_enq_valid = auto_out_d_valid & _T_395; 
  assign Queue_1_io_enq_bits_id = auto_out_d_bits_source[2:2]; 
  assign Queue_1_io_enq_bits_resp = _T_371 ? 2'h2 : 2'h0; 
  assign Queue_1_io_deq_ready = auto_in_bready & _T_403; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_54_0 = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_54_1 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_260 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_270 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_325_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_209_0 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_209_1 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_325_1 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_382 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_402_0 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_402_1 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_54_0 <= 2'h0;
    end else begin
      if (_T_150) begin
        _T_54_0 <= _T_152;
      end
    end
    if (reset) begin
      _T_54_1 <= 2'h0;
    end else begin
      if (_T_154) begin
        _T_54_1 <= _T_156;
      end
    end
    if (reset) begin
      _T_260 <= 8'h0;
    end else begin
      if (_T_262) begin
        if (_T_296) begin
          _T_260 <= auto_in_awlen;
        end else begin
          _T_260 <= 8'h0;
        end
      end else begin
        _T_260 <= _T_322;
      end
    end
    if (reset) begin
      _T_270 <= 2'h3;
    end else begin
      if (_T_285) begin
        _T_270 <= _T_289;
      end
    end
    if (reset) begin
      _T_325_0 <= 1'h0;
    end else begin
      if (_T_261) begin
        _T_325_0 <= _T_295;
      end
    end
    if (reset) begin
      _T_209_0 <= 2'h0;
    end else begin
      if (_T_253) begin
        _T_209_0 <= _T_255;
      end
    end
    if (reset) begin
      _T_209_1 <= 2'h0;
    end else begin
      if (_T_257) begin
        _T_209_1 <= _T_259;
      end
    end
    if (reset) begin
      _T_325_1 <= 1'h0;
    end else begin
      if (_T_261) begin
        _T_325_1 <= _T_296;
      end
    end
    if (reset) begin
      _T_382 <= 3'h0;
    end else begin
      if (_T_374) begin
        if (_T_385) begin
          if (_T_373) begin
            _T_382 <= _T_379;
          end else begin
            _T_382 <= 3'h0;
          end
        end else begin
          _T_382 <= _T_384;
        end
      end
    end
    if (reset) begin
      _T_402_0 <= 2'h0;
    end else begin
      if (_T_410) begin
        _T_402_0 <= _T_412;
      end
    end
    if (reset) begin
      _T_402_1 <= 2'h0;
    end else begin
      if (_T_414) begin
        _T_402_1 <= _T_416;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_67) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToTL.scala:88 assert (!in.ar.valid || r_size1 === UIntToOH1(r_size, beatCountBits)) // because aligned\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_67) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_222) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToTL.scala:107 assert (!in.aw.valid || w_size1 === UIntToOH1(w_size, beatCountBits)) // because aligned\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_222) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_230) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToTL.scala:108 assert (!in.aw.valid || in.aw.bits.len === UInt(0) || in.aw.bits.size === UInt(log2Ceil(beatBytes))) // because aligned\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_230) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_268) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_268) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_309) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_309) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_316) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:70 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_316) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_AXI4UserYanker_1( 
  input         clock, 
  input         reset, 
  output        auto_in_awready, 
  input         auto_in_awvalid, 
  input  [30:0] auto_in_awaddr, 
  input  [7:0]  auto_in_awlen, 
  input  [2:0]  auto_in_awsize, 
  input  [1:0]  auto_in_awburst, 
  input         auto_in_awlock, 
  input  [3:0]  auto_in_awcache, 
  input  [2:0]  auto_in_awprot, 
  input  [3:0]  auto_in_awqos, 
  input  [15:0] auto_in_awuser, 
  input  [63:0] auto_in_awinstret, 
  output        auto_in_wready, 
  input         auto_in_wvalid, 
  input  [63:0] auto_in_wdata, 
  input  [7:0]  auto_in_wstrb, 
  input         auto_in_wlast, 
  input         auto_in_bready, 
  output        auto_in_bvalid, 
  output [1:0]  auto_in_bresp, 
  output [15:0] auto_in_buser, 
  output        auto_in_arready, 
  input         auto_in_arvalid, 
  input  [30:0] auto_in_araddr, 
  input  [7:0]  auto_in_arlen, 
  input  [2:0]  auto_in_arsize, 
  input  [1:0]  auto_in_arburst, 
  input         auto_in_arlock, 
  input  [3:0]  auto_in_arcache, 
  input  [2:0]  auto_in_arprot, 
  input  [3:0]  auto_in_arqos, 
  input  [15:0] auto_in_aruser, 
  input  [63:0] auto_in_arinstret, 
  input         auto_in_rready, 
  output        auto_in_rvalid, 
  output [63:0] auto_in_rdata, 
  output [1:0]  auto_in_rresp, 
  output [15:0] auto_in_ruser, 
  output        auto_in_rlast, 
  input         auto_out_awready, 
  output        auto_out_awvalid, 
  output [30:0] auto_out_awaddr, 
  output [7:0]  auto_out_awlen, 
  output [2:0]  auto_out_awsize, 
  output [1:0]  auto_out_awburst, 
  output        auto_out_awlock, 
  output [3:0]  auto_out_awcache, 
  output [2:0]  auto_out_awprot, 
  output [3:0]  auto_out_awqos, 
  output [63:0] auto_out_awinstret, 
  input         auto_out_wready, 
  output        auto_out_wvalid, 
  output [63:0] auto_out_wdata, 
  output [7:0]  auto_out_wstrb, 
  output        auto_out_wlast, 
  output        auto_out_bready, 
  input         auto_out_bvalid, 
  input  [1:0]  auto_out_bresp, 
  input         auto_out_arready, 
  output        auto_out_arvalid, 
  output [30:0] auto_out_araddr, 
  output [7:0]  auto_out_arlen, 
  output [2:0]  auto_out_arsize, 
  output [1:0]  auto_out_arburst, 
  output        auto_out_arlock, 
  output [3:0]  auto_out_arcache, 
  output [2:0]  auto_out_arprot, 
  output [3:0]  auto_out_arqos, 
  output [63:0] auto_out_arinstret, 
  output        auto_out_rready, 
  input         auto_out_rvalid, 
  input  [63:0] auto_out_rdata, 
  input  [1:0]  auto_out_rresp, 
  input         auto_out_rlast 
);
  wire  Queue_clock; 
  wire  Queue_reset; 
  wire  Queue_io_enq_ready; 
  wire  Queue_io_enq_valid; 
  wire [15:0] Queue_io_enq_bits; 
  wire  Queue_io_deq_ready; 
  wire  Queue_io_deq_valid; 
  wire [15:0] Queue_io_deq_bits; 
  wire  Queue_1_clock; 
  wire  Queue_1_reset; 
  wire  Queue_1_io_enq_ready; 
  wire  Queue_1_io_enq_valid; 
  wire [15:0] Queue_1_io_enq_bits; 
  wire  Queue_1_io_deq_ready; 
  wire  Queue_1_io_deq_valid; 
  wire [15:0] Queue_1_io_deq_bits; 
  wire  _T_2_0; 
  wire  _T_7; 
  wire  _T_5_0; 
  wire  _T_8; 
  wire  _T_10; 
  wire  _T_11; 
  wire  _T_12; 
  wire  _T_17_0; 
  wire  _T_22; 
  wire  _T_20_0; 
  wire  _T_23; 
  wire  _T_25; 
  wire  _T_26; 
  dual_Queue_53 dual_Queue ( 
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits(Queue_io_enq_bits),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits(Queue_io_deq_bits)
  );
  dual_Queue_53 Queue_1 ( 
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits(Queue_1_io_enq_bits),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits(Queue_1_io_deq_bits)
  );
  assign _T_2_0 = Queue_io_enq_ready; 
  assign _T_7 = auto_out_rvalid == 1'h0; 
  assign _T_5_0 = Queue_io_deq_valid; 
  assign _T_8 = _T_7 | _T_5_0; 
  assign _T_10 = _T_8 | reset; 
  assign _T_11 = _T_10 == 1'h0; 
  assign _T_12 = auto_out_rvalid & auto_in_rready; 
  assign _T_17_0 = Queue_1_io_enq_ready; 
  assign _T_22 = auto_out_bvalid == 1'h0; 
  assign _T_20_0 = Queue_1_io_deq_valid; 
  assign _T_23 = _T_22 | _T_20_0; 
  assign _T_25 = _T_23 | reset; 
  assign _T_26 = _T_25 == 1'h0; 
  assign auto_in_awready = auto_out_awready & _T_17_0; 
  assign auto_in_wready = auto_out_wready; 
  assign auto_in_bvalid = auto_out_bvalid; 
  assign auto_in_bresp = auto_out_bresp; 
  assign auto_in_buser = Queue_1_io_deq_bits; 
  assign auto_in_arready = auto_out_arready & _T_2_0; 
  assign auto_in_rvalid = auto_out_rvalid; 
  assign auto_in_rdata = auto_out_rdata; 
  assign auto_in_rresp = auto_out_rresp; 
  assign auto_in_ruser = Queue_io_deq_bits; 
  assign auto_in_rlast = auto_out_rlast; 
  assign auto_out_awvalid = auto_in_awvalid & _T_17_0; 
  assign auto_out_awaddr = auto_in_awaddr; 
  assign auto_out_awlen = auto_in_awlen; 
  assign auto_out_awsize = auto_in_awsize; 
  assign auto_out_awburst = auto_in_awburst; 
  assign auto_out_awlock = auto_in_awlock; 
  assign auto_out_awcache = auto_in_awcache; 
  assign auto_out_awprot = auto_in_awprot; 
  assign auto_out_awqos = auto_in_awqos; 
  assign auto_out_awinstret = auto_in_awinstret; 
  assign auto_out_wvalid = auto_in_wvalid; 
  assign auto_out_wdata = auto_in_wdata; 
  assign auto_out_wstrb = auto_in_wstrb; 
  assign auto_out_wlast = auto_in_wlast; 
  assign auto_out_bready = auto_in_bready; 
  assign auto_out_arvalid = auto_in_arvalid & _T_2_0; 
  assign auto_out_araddr = auto_in_araddr; 
  assign auto_out_arlen = auto_in_arlen; 
  assign auto_out_arsize = auto_in_arsize; 
  assign auto_out_arburst = auto_in_arburst; 
  assign auto_out_arlock = auto_in_arlock; 
  assign auto_out_arcache = auto_in_arcache; 
  assign auto_out_arprot = auto_in_arprot; 
  assign auto_out_arqos = auto_in_arqos; 
  assign auto_out_arinstret = auto_in_arinstret; 
  assign auto_out_rready = auto_in_rready; 
  assign Queue_clock = clock; 
  assign Queue_reset = reset; 
  assign Queue_io_enq_valid = auto_in_arvalid & auto_out_arready; 
  assign Queue_io_enq_bits = auto_in_aruser; 
  assign Queue_io_deq_ready = _T_12 & auto_out_rlast; 
  assign Queue_1_clock = clock; 
  assign Queue_1_reset = reset; 
  assign Queue_1_io_enq_valid = auto_in_awvalid & auto_out_awready; 
  assign Queue_1_io_enq_bits = auto_in_awuser; 
  assign Queue_1_io_deq_ready = auto_out_bvalid & auto_in_bready; 
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_11) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:54 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_11) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_26) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:75 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_26) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_AXI4UserYanker_2( 
  input         clock, 
  input         reset, 
  output        auto_in_awready, 
  input         auto_in_awvalid, 
  input         auto_in_awid, 
  input  [31:0] auto_in_awaddr, 
  input  [7:0]  auto_in_awlen, 
  input  [2:0]  auto_in_awsize, 
  input  [16:0] auto_in_awuser, 
  output        auto_in_wready, 
  input         auto_in_wvalid, 
  input  [63:0] auto_in_wdata, 
  input  [7:0]  auto_in_wstrb, 
  input         auto_in_wlast, 
  input         auto_in_bready, 
  output        auto_in_bvalid, 
  output        auto_in_bid, 
  output [1:0]  auto_in_bresp, 
  output [16:0] auto_in_buser, 
  output        auto_in_arready, 
  input         auto_in_arvalid, 
  input         auto_in_arid, 
  input  [31:0] auto_in_araddr, 
  input  [7:0]  auto_in_arlen, 
  input  [2:0]  auto_in_arsize, 
  input  [16:0] auto_in_aruser, 
  input         auto_in_rready, 
  output        auto_in_rvalid, 
  output        auto_in_rid, 
  output [63:0] auto_in_rdata, 
  output [1:0]  auto_in_rresp, 
  output [16:0] auto_in_ruser, 
  output        auto_in_rlast, 
  input         auto_out_awready, 
  output        auto_out_awvalid, 
  output        auto_out_awid, 
  output [31:0] auto_out_awaddr, 
  output [7:0]  auto_out_awlen, 
  output [2:0]  auto_out_awsize, 
  input         auto_out_wready, 
  output        auto_out_wvalid, 
  output [63:0] auto_out_wdata, 
  output [7:0]  auto_out_wstrb, 
  output        auto_out_wlast, 
  output        auto_out_bready, 
  input         auto_out_bvalid, 
  input         auto_out_bid, 
  input  [1:0]  auto_out_bresp, 
  input         auto_out_arready, 
  output        auto_out_arvalid, 
  output        auto_out_arid, 
  output [31:0] auto_out_araddr, 
  output [7:0]  auto_out_arlen, 
  output [2:0]  auto_out_arsize, 
  output        auto_out_rready, 
  input         auto_out_rvalid, 
  input         auto_out_rid, 
  input  [63:0] auto_out_rdata, 
  input  [1:0]  auto_out_rresp, 
  input         auto_out_rlast 
);
  wire  Queue_clock; 
  wire  Queue_reset; 
  wire  Queue_io_enq_ready; 
  wire  Queue_io_enq_valid; 
  wire [16:0] Queue_io_enq_bits; 
  wire  Queue_io_deq_ready; 
  wire  Queue_io_deq_valid; 
  wire [16:0] Queue_io_deq_bits; 
  wire  Queue_1_clock; 
  wire  Queue_1_reset; 
  wire  Queue_1_io_enq_ready; 
  wire  Queue_1_io_enq_valid; 
  wire [16:0] Queue_1_io_enq_bits; 
  wire  Queue_1_io_deq_ready; 
  wire  Queue_1_io_deq_valid; 
  wire [16:0] Queue_1_io_deq_bits; 
  wire  Queue_2_clock; 
  wire  Queue_2_reset; 
  wire  Queue_2_io_enq_ready; 
  wire  Queue_2_io_enq_valid; 
  wire [16:0] Queue_2_io_enq_bits; 
  wire  Queue_2_io_deq_ready; 
  wire  Queue_2_io_deq_valid; 
  wire [16:0] Queue_2_io_deq_bits; 
  wire  Queue_3_clock; 
  wire  Queue_3_reset; 
  wire  Queue_3_io_enq_ready; 
  wire  Queue_3_io_enq_valid; 
  wire [16:0] Queue_3_io_enq_bits; 
  wire  Queue_3_io_deq_ready; 
  wire  Queue_3_io_deq_valid; 
  wire [16:0] Queue_3_io_deq_bits; 
  wire  _T_2_0; 
  wire  _T_2_1; 
  wire  _GEN_1; 
  wire  _T_7; 
  wire  _T_5_0; 
  wire  _T_5_1; 
  wire  _GEN_3; 
  wire  _T_8; 
  wire  _T_10; 
  wire  _T_11; 
  wire [16:0] _T_6_0; 
  wire [16:0] _T_6_1; 
  wire [1:0] _T_13; 
  wire  _T_15; 
  wire  _T_16; 
  wire [1:0] _T_18; 
  wire  _T_20; 
  wire  _T_21; 
  wire  _T_22; 
  wire  _T_23; 
  wire  _T_25; 
  wire  _T_28; 
  wire  _T_32_0; 
  wire  _T_32_1; 
  wire  _GEN_7; 
  wire  _T_37; 
  wire  _T_35_0; 
  wire  _T_35_1; 
  wire  _GEN_9; 
  wire  _T_38; 
  wire  _T_40; 
  wire  _T_41; 
  wire [16:0] _T_36_0; 
  wire [16:0] _T_36_1; 
  wire [1:0] _T_43; 
  wire  _T_45; 
  wire  _T_46; 
  wire [1:0] _T_48; 
  wire  _T_50; 
  wire  _T_51; 
  wire  _T_52; 
  wire  _T_54; 
  dual_Queue_60 dual_Queue ( 
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits(Queue_io_enq_bits),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits(Queue_io_deq_bits)
  );
  dual_Queue_60 Queue_1 ( 
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits(Queue_1_io_enq_bits),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits(Queue_1_io_deq_bits)
  );
  dual_Queue_60 dual_Queue_2 ( 
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits(Queue_2_io_enq_bits),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits(Queue_2_io_deq_bits)
  );
  dual_Queue_60 Queue_3 ( 
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits(Queue_3_io_enq_bits),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits(Queue_3_io_deq_bits)
  );
  assign _T_2_0 = Queue_io_enq_ready; 
  assign _T_2_1 = Queue_1_io_enq_ready; 
  assign _GEN_1 = auto_in_arid ? _T_2_1 : _T_2_0; 
  assign _T_7 = auto_out_rvalid == 1'h0; 
  assign _T_5_0 = Queue_io_deq_valid; 
  assign _T_5_1 = Queue_1_io_deq_valid; 
  assign _GEN_3 = auto_out_rid ? _T_5_1 : _T_5_0; 
  assign _T_8 = _T_7 | _GEN_3; 
  assign _T_10 = _T_8 | reset; 
  assign _T_11 = _T_10 == 1'h0; 
  assign _T_6_0 = Queue_io_deq_bits; 
  assign _T_6_1 = Queue_1_io_deq_bits; 
  assign _T_13 = 2'h1 << auto_in_arid; 
  assign _T_15 = _T_13[0]; 
  assign _T_16 = _T_13[1]; 
  assign _T_18 = 2'h1 << auto_out_rid; 
  assign _T_20 = _T_18[0]; 
  assign _T_21 = _T_18[1]; 
  assign _T_22 = auto_out_rvalid & auto_in_rready; 
  assign _T_23 = _T_22 & _T_20; 
  assign _T_25 = auto_in_arvalid & auto_out_arready; 
  assign _T_28 = _T_22 & _T_21; 
  assign _T_32_0 = Queue_2_io_enq_ready; 
  assign _T_32_1 = Queue_3_io_enq_ready; 
  assign _GEN_7 = auto_in_awid ? _T_32_1 : _T_32_0; 
  assign _T_37 = auto_out_bvalid == 1'h0; 
  assign _T_35_0 = Queue_2_io_deq_valid; 
  assign _T_35_1 = Queue_3_io_deq_valid; 
  assign _GEN_9 = auto_out_bid ? _T_35_1 : _T_35_0; 
  assign _T_38 = _T_37 | _GEN_9; 
  assign _T_40 = _T_38 | reset; 
  assign _T_41 = _T_40 == 1'h0; 
  assign _T_36_0 = Queue_2_io_deq_bits; 
  assign _T_36_1 = Queue_3_io_deq_bits; 
  assign _T_43 = 2'h1 << auto_in_awid; 
  assign _T_45 = _T_43[0]; 
  assign _T_46 = _T_43[1]; 
  assign _T_48 = 2'h1 << auto_out_bid; 
  assign _T_50 = _T_48[0]; 
  assign _T_51 = _T_48[1]; 
  assign _T_52 = auto_out_bvalid & auto_in_bready; 
  assign _T_54 = auto_in_awvalid & auto_out_awready; 
  assign auto_in_awready = auto_out_awready & _GEN_7; 
  assign auto_in_wready = auto_out_wready; 
  assign auto_in_bvalid = auto_out_bvalid; 
  assign auto_in_bid = auto_out_bid; 
  assign auto_in_bresp = auto_out_bresp; 
  assign auto_in_buser = auto_out_bid ? _T_36_1 : _T_36_0; 
  assign auto_in_arready = auto_out_arready & _GEN_1; 
  assign auto_in_rvalid = auto_out_rvalid; 
  assign auto_in_rid = auto_out_rid; 
  assign auto_in_rdata = auto_out_rdata; 
  assign auto_in_rresp = auto_out_rresp; 
  assign auto_in_ruser = auto_out_rid ? _T_6_1 : _T_6_0; 
  assign auto_in_rlast = auto_out_rlast; 
  assign auto_out_awvalid = auto_in_awvalid & _GEN_7; 
  assign auto_out_awid = auto_in_awid; 
  assign auto_out_awaddr = auto_in_awaddr; 
  assign auto_out_awlen = auto_in_awlen; 
  assign auto_out_awsize = auto_in_awsize; 
  assign auto_out_wvalid = auto_in_wvalid; 
  assign auto_out_wdata = auto_in_wdata; 
  assign auto_out_wstrb = auto_in_wstrb; 
  assign auto_out_wlast = auto_in_wlast; 
  assign auto_out_bready = auto_in_bready; 
  assign auto_out_arvalid = auto_in_arvalid & _GEN_1; 
  assign auto_out_arid = auto_in_arid; 
  assign auto_out_araddr = auto_in_araddr; 
  assign auto_out_arlen = auto_in_arlen; 
  assign auto_out_arsize = auto_in_arsize; 
  assign auto_out_rready = auto_in_rready; 
  assign Queue_clock = clock; 
  assign Queue_reset = reset; 
  assign Queue_io_enq_valid = _T_25 & _T_15; 
  assign Queue_io_enq_bits = auto_in_aruser; 
  assign Queue_io_deq_ready = _T_23 & auto_out_rlast; 
  assign Queue_1_clock = clock; 
  assign Queue_1_reset = reset; 
  assign Queue_1_io_enq_valid = _T_25 & _T_16; 
  assign Queue_1_io_enq_bits = auto_in_aruser; 
  assign Queue_1_io_deq_ready = _T_28 & auto_out_rlast; 
  assign Queue_2_clock = clock; 
  assign Queue_2_reset = reset; 
  assign Queue_2_io_enq_valid = _T_54 & _T_45; 
  assign Queue_2_io_enq_bits = auto_in_awuser; 
  assign Queue_2_io_deq_ready = _T_52 & _T_50; 
  assign Queue_3_clock = clock; 
  assign Queue_3_reset = reset; 
  assign Queue_3_io_enq_valid = _T_54 & _T_46; 
  assign Queue_3_io_enq_bits = auto_in_awuser; 
  assign Queue_3_io_deq_ready = _T_52 & _T_51; 
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_11) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:54 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_11) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_41) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:75 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_41) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_AXI4UserYanker( 
  input         clock, 
  input         reset, 
  output        auto_in_awready, 
  input         auto_in_awvalid, 
  input  [3:0]  auto_in_awid, 
  input  [31:0] auto_in_awaddr, 
  input  [7:0]  auto_in_awlen, 
  input  [2:0]  auto_in_awsize, 
  input  [1:0]  auto_in_awburst, 
  input         auto_in_awlock, 
  input  [3:0]  auto_in_awcache, 
  input  [2:0]  auto_in_awprot, 
  input  [3:0]  auto_in_awqos, 
  input  [11:0] auto_in_awuser, 
  input  [63:0] auto_in_awinstret, 
  output        auto_in_wready, 
  input         auto_in_wvalid, 
  input  [63:0] auto_in_wdata, 
  input  [7:0]  auto_in_wstrb, 
  input         auto_in_wlast, 
  input         auto_in_bready, 
  output        auto_in_bvalid, 
  output [3:0]  auto_in_bid, 
  output [1:0]  auto_in_bresp, 
  output [11:0] auto_in_buser, 
  output        auto_in_arready, 
  input         auto_in_arvalid, 
  input  [3:0]  auto_in_arid, 
  input  [31:0] auto_in_araddr, 
  input  [7:0]  auto_in_arlen, 
  input  [2:0]  auto_in_arsize, 
  input  [1:0]  auto_in_arburst, 
  input         auto_in_arlock, 
  input  [3:0]  auto_in_arcache, 
  input  [2:0]  auto_in_arprot, 
  input  [3:0]  auto_in_arqos, 
  input  [11:0] auto_in_aruser, 
  input  [63:0] auto_in_arinstret, 
  input         auto_in_rready, 
  output        auto_in_rvalid, 
  output [3:0]  auto_in_rid, 
  output [63:0] auto_in_rdata, 
  output [1:0]  auto_in_rresp, 
  output [11:0] auto_in_ruser, 
  output        auto_in_rlast, 
  input         auto_out_awready, 
  output        auto_out_awvalid, 
  output [3:0]  auto_out_awid, 
  output [31:0] auto_out_awaddr, 
  output [7:0]  auto_out_awlen, 
  output [2:0]  auto_out_awsize, 
  output [1:0]  auto_out_awburst, 
  output        auto_out_awlock, 
  output [3:0]  auto_out_awcache, 
  output [2:0]  auto_out_awprot, 
  output [3:0]  auto_out_awqos, 
  output [63:0] auto_out_awinstret, 
  input         auto_out_wready, 
  output        auto_out_wvalid, 
  output [63:0] auto_out_wdata, 
  output [7:0]  auto_out_wstrb, 
  output        auto_out_wlast, 
  output        auto_out_bready, 
  input         auto_out_bvalid, 
  input  [3:0]  auto_out_bid, 
  input  [1:0]  auto_out_bresp, 
  input         auto_out_arready, 
  output        auto_out_arvalid, 
  output [3:0]  auto_out_arid, 
  output [31:0] auto_out_araddr, 
  output [7:0]  auto_out_arlen, 
  output [2:0]  auto_out_arsize, 
  output [1:0]  auto_out_arburst, 
  output        auto_out_arlock, 
  output [3:0]  auto_out_arcache, 
  output [2:0]  auto_out_arprot, 
  output [3:0]  auto_out_arqos, 
  output [63:0] auto_out_arinstret, 
  output        auto_out_rready, 
  input         auto_out_rvalid, 
  input  [3:0]  auto_out_rid, 
  input  [63:0] auto_out_rdata, 
  input  [1:0]  auto_out_rresp, 
  input         auto_out_rlast 
);
  wire  Queue_clock; 
  wire  Queue_reset; 
  wire  Queue_io_enq_ready; 
  wire  Queue_io_enq_valid; 
  wire [11:0] Queue_io_enq_bits; 
  wire  Queue_io_deq_ready; 
  wire  Queue_io_deq_valid; 
  wire [11:0] Queue_io_deq_bits; 
  wire  Queue_1_clock; 
  wire  Queue_1_reset; 
  wire  Queue_1_io_enq_ready; 
  wire  Queue_1_io_enq_valid; 
  wire [11:0] Queue_1_io_enq_bits; 
  wire  Queue_1_io_deq_ready; 
  wire  Queue_1_io_deq_valid; 
  wire [11:0] Queue_1_io_deq_bits; 
  wire  Queue_2_clock; 
  wire  Queue_2_reset; 
  wire  Queue_2_io_enq_ready; 
  wire  Queue_2_io_enq_valid; 
  wire [11:0] Queue_2_io_enq_bits; 
  wire  Queue_2_io_deq_ready; 
  wire  Queue_2_io_deq_valid; 
  wire [11:0] Queue_2_io_deq_bits; 
  wire  Queue_3_clock; 
  wire  Queue_3_reset; 
  wire  Queue_3_io_enq_ready; 
  wire  Queue_3_io_enq_valid; 
  wire [11:0] Queue_3_io_enq_bits; 
  wire  Queue_3_io_deq_ready; 
  wire  Queue_3_io_deq_valid; 
  wire [11:0] Queue_3_io_deq_bits; 
  wire  Queue_4_clock; 
  wire  Queue_4_reset; 
  wire  Queue_4_io_enq_ready; 
  wire  Queue_4_io_enq_valid; 
  wire [11:0] Queue_4_io_enq_bits; 
  wire  Queue_4_io_deq_ready; 
  wire  Queue_4_io_deq_valid; 
  wire [11:0] Queue_4_io_deq_bits; 
  wire  Queue_5_clock; 
  wire  Queue_5_reset; 
  wire  Queue_5_io_enq_ready; 
  wire  Queue_5_io_enq_valid; 
  wire [11:0] Queue_5_io_enq_bits; 
  wire  Queue_5_io_deq_ready; 
  wire  Queue_5_io_deq_valid; 
  wire [11:0] Queue_5_io_deq_bits; 
  wire  Queue_6_clock; 
  wire  Queue_6_reset; 
  wire  Queue_6_io_enq_ready; 
  wire  Queue_6_io_enq_valid; 
  wire [11:0] Queue_6_io_enq_bits; 
  wire  Queue_6_io_deq_ready; 
  wire  Queue_6_io_deq_valid; 
  wire [11:0] Queue_6_io_deq_bits; 
  wire  Queue_7_clock; 
  wire  Queue_7_reset; 
  wire  Queue_7_io_enq_ready; 
  wire  Queue_7_io_enq_valid; 
  wire [11:0] Queue_7_io_enq_bits; 
  wire  Queue_7_io_deq_ready; 
  wire  Queue_7_io_deq_valid; 
  wire [11:0] Queue_7_io_deq_bits; 
  wire  Queue_8_clock; 
  wire  Queue_8_reset; 
  wire  Queue_8_io_enq_ready; 
  wire  Queue_8_io_enq_valid; 
  wire [11:0] Queue_8_io_enq_bits; 
  wire  Queue_8_io_deq_ready; 
  wire  Queue_8_io_deq_valid; 
  wire [11:0] Queue_8_io_deq_bits; 
  wire  Queue_9_clock; 
  wire  Queue_9_reset; 
  wire  Queue_9_io_enq_ready; 
  wire  Queue_9_io_enq_valid; 
  wire [11:0] Queue_9_io_enq_bits; 
  wire  Queue_9_io_deq_ready; 
  wire  Queue_9_io_deq_valid; 
  wire [11:0] Queue_9_io_deq_bits; 
  wire  Queue_10_clock; 
  wire  Queue_10_reset; 
  wire  Queue_10_io_enq_ready; 
  wire  Queue_10_io_enq_valid; 
  wire [11:0] Queue_10_io_enq_bits; 
  wire  Queue_10_io_deq_ready; 
  wire  Queue_10_io_deq_valid; 
  wire [11:0] Queue_10_io_deq_bits; 
  wire  Queue_11_clock; 
  wire  Queue_11_reset; 
  wire  Queue_11_io_enq_ready; 
  wire  Queue_11_io_enq_valid; 
  wire [11:0] Queue_11_io_enq_bits; 
  wire  Queue_11_io_deq_ready; 
  wire  Queue_11_io_deq_valid; 
  wire [11:0] Queue_11_io_deq_bits; 
  wire  Queue_12_clock; 
  wire  Queue_12_reset; 
  wire  Queue_12_io_enq_ready; 
  wire  Queue_12_io_enq_valid; 
  wire [11:0] Queue_12_io_enq_bits; 
  wire  Queue_12_io_deq_ready; 
  wire  Queue_12_io_deq_valid; 
  wire [11:0] Queue_12_io_deq_bits; 
  wire  Queue_13_clock; 
  wire  Queue_13_reset; 
  wire  Queue_13_io_enq_ready; 
  wire  Queue_13_io_enq_valid; 
  wire [11:0] Queue_13_io_enq_bits; 
  wire  Queue_13_io_deq_ready; 
  wire  Queue_13_io_deq_valid; 
  wire [11:0] Queue_13_io_deq_bits; 
  wire  Queue_14_clock; 
  wire  Queue_14_reset; 
  wire  Queue_14_io_enq_ready; 
  wire  Queue_14_io_enq_valid; 
  wire [11:0] Queue_14_io_enq_bits; 
  wire  Queue_14_io_deq_ready; 
  wire  Queue_14_io_deq_valid; 
  wire [11:0] Queue_14_io_deq_bits; 
  wire  Queue_15_clock; 
  wire  Queue_15_reset; 
  wire  Queue_15_io_enq_ready; 
  wire  Queue_15_io_enq_valid; 
  wire [11:0] Queue_15_io_enq_bits; 
  wire  Queue_15_io_deq_ready; 
  wire  Queue_15_io_deq_valid; 
  wire [11:0] Queue_15_io_deq_bits; 
  wire  Queue_16_clock; 
  wire  Queue_16_reset; 
  wire  Queue_16_io_enq_ready; 
  wire  Queue_16_io_enq_valid; 
  wire [11:0] Queue_16_io_enq_bits; 
  wire  Queue_16_io_deq_ready; 
  wire  Queue_16_io_deq_valid; 
  wire [11:0] Queue_16_io_deq_bits; 
  wire  Queue_17_clock; 
  wire  Queue_17_reset; 
  wire  Queue_17_io_enq_ready; 
  wire  Queue_17_io_enq_valid; 
  wire [11:0] Queue_17_io_enq_bits; 
  wire  Queue_17_io_deq_ready; 
  wire  Queue_17_io_deq_valid; 
  wire [11:0] Queue_17_io_deq_bits; 
  wire  Queue_18_clock; 
  wire  Queue_18_reset; 
  wire  Queue_18_io_enq_ready; 
  wire  Queue_18_io_enq_valid; 
  wire [11:0] Queue_18_io_enq_bits; 
  wire  Queue_18_io_deq_ready; 
  wire  Queue_18_io_deq_valid; 
  wire [11:0] Queue_18_io_deq_bits; 
  wire  Queue_19_clock; 
  wire  Queue_19_reset; 
  wire  Queue_19_io_enq_ready; 
  wire  Queue_19_io_enq_valid; 
  wire [11:0] Queue_19_io_enq_bits; 
  wire  Queue_19_io_deq_ready; 
  wire  Queue_19_io_deq_valid; 
  wire [11:0] Queue_19_io_deq_bits; 
  wire  Queue_20_clock; 
  wire  Queue_20_reset; 
  wire  Queue_20_io_enq_ready; 
  wire  Queue_20_io_enq_valid; 
  wire [11:0] Queue_20_io_enq_bits; 
  wire  Queue_20_io_deq_ready; 
  wire  Queue_20_io_deq_valid; 
  wire [11:0] Queue_20_io_deq_bits; 
  wire  Queue_21_clock; 
  wire  Queue_21_reset; 
  wire  Queue_21_io_enq_ready; 
  wire  Queue_21_io_enq_valid; 
  wire [11:0] Queue_21_io_enq_bits; 
  wire  Queue_21_io_deq_ready; 
  wire  Queue_21_io_deq_valid; 
  wire [11:0] Queue_21_io_deq_bits; 
  wire  Queue_22_clock; 
  wire  Queue_22_reset; 
  wire  Queue_22_io_enq_ready; 
  wire  Queue_22_io_enq_valid; 
  wire [11:0] Queue_22_io_enq_bits; 
  wire  Queue_22_io_deq_ready; 
  wire  Queue_22_io_deq_valid; 
  wire [11:0] Queue_22_io_deq_bits; 
  wire  Queue_23_clock; 
  wire  Queue_23_reset; 
  wire  Queue_23_io_enq_ready; 
  wire  Queue_23_io_enq_valid; 
  wire [11:0] Queue_23_io_enq_bits; 
  wire  Queue_23_io_deq_ready; 
  wire  Queue_23_io_deq_valid; 
  wire [11:0] Queue_23_io_deq_bits; 
  wire  Queue_24_clock; 
  wire  Queue_24_reset; 
  wire  Queue_24_io_enq_ready; 
  wire  Queue_24_io_enq_valid; 
  wire [11:0] Queue_24_io_enq_bits; 
  wire  Queue_24_io_deq_ready; 
  wire  Queue_24_io_deq_valid; 
  wire [11:0] Queue_24_io_deq_bits; 
  wire  Queue_25_clock; 
  wire  Queue_25_reset; 
  wire  Queue_25_io_enq_ready; 
  wire  Queue_25_io_enq_valid; 
  wire [11:0] Queue_25_io_enq_bits; 
  wire  Queue_25_io_deq_ready; 
  wire  Queue_25_io_deq_valid; 
  wire [11:0] Queue_25_io_deq_bits; 
  wire  Queue_26_clock; 
  wire  Queue_26_reset; 
  wire  Queue_26_io_enq_ready; 
  wire  Queue_26_io_enq_valid; 
  wire [11:0] Queue_26_io_enq_bits; 
  wire  Queue_26_io_deq_ready; 
  wire  Queue_26_io_deq_valid; 
  wire [11:0] Queue_26_io_deq_bits; 
  wire  Queue_27_clock; 
  wire  Queue_27_reset; 
  wire  Queue_27_io_enq_ready; 
  wire  Queue_27_io_enq_valid; 
  wire [11:0] Queue_27_io_enq_bits; 
  wire  Queue_27_io_deq_ready; 
  wire  Queue_27_io_deq_valid; 
  wire [11:0] Queue_27_io_deq_bits; 
  wire  Queue_28_clock; 
  wire  Queue_28_reset; 
  wire  Queue_28_io_enq_ready; 
  wire  Queue_28_io_enq_valid; 
  wire [11:0] Queue_28_io_enq_bits; 
  wire  Queue_28_io_deq_ready; 
  wire  Queue_28_io_deq_valid; 
  wire [11:0] Queue_28_io_deq_bits; 
  wire  Queue_29_clock; 
  wire  Queue_29_reset; 
  wire  Queue_29_io_enq_ready; 
  wire  Queue_29_io_enq_valid; 
  wire [11:0] Queue_29_io_enq_bits; 
  wire  Queue_29_io_deq_ready; 
  wire  Queue_29_io_deq_valid; 
  wire [11:0] Queue_29_io_deq_bits; 
  wire  Queue_30_clock; 
  wire  Queue_30_reset; 
  wire  Queue_30_io_enq_ready; 
  wire  Queue_30_io_enq_valid; 
  wire [11:0] Queue_30_io_enq_bits; 
  wire  Queue_30_io_deq_ready; 
  wire  Queue_30_io_deq_valid; 
  wire [11:0] Queue_30_io_deq_bits; 
  wire  Queue_31_clock; 
  wire  Queue_31_reset; 
  wire  Queue_31_io_enq_ready; 
  wire  Queue_31_io_enq_valid; 
  wire [11:0] Queue_31_io_enq_bits; 
  wire  Queue_31_io_deq_ready; 
  wire  Queue_31_io_deq_valid; 
  wire [11:0] Queue_31_io_deq_bits; 
  wire  _T_2_0; 
  wire  _T_2_1; 
  wire  _GEN_1; 
  wire  _T_2_2; 
  wire  _GEN_2; 
  wire  _T_2_3; 
  wire  _GEN_3; 
  wire  _T_2_4; 
  wire  _GEN_4; 
  wire  _T_2_5; 
  wire  _GEN_5; 
  wire  _T_2_6; 
  wire  _GEN_6; 
  wire  _T_2_7; 
  wire  _GEN_7; 
  wire  _T_2_8; 
  wire  _GEN_8; 
  wire  _T_2_9; 
  wire  _GEN_9; 
  wire  _T_2_10; 
  wire  _GEN_10; 
  wire  _T_2_11; 
  wire  _GEN_11; 
  wire  _T_2_12; 
  wire  _GEN_12; 
  wire  _T_2_13; 
  wire  _GEN_13; 
  wire  _T_2_14; 
  wire  _GEN_14; 
  wire  _T_2_15; 
  wire  _GEN_15; 
  wire  _T_7; 
  wire  _T_5_0; 
  wire  _T_5_1; 
  wire  _GEN_17; 
  wire  _T_5_2; 
  wire  _GEN_18; 
  wire  _T_5_3; 
  wire  _GEN_19; 
  wire  _T_5_4; 
  wire  _GEN_20; 
  wire  _T_5_5; 
  wire  _GEN_21; 
  wire  _T_5_6; 
  wire  _GEN_22; 
  wire  _T_5_7; 
  wire  _GEN_23; 
  wire  _T_5_8; 
  wire  _GEN_24; 
  wire  _T_5_9; 
  wire  _GEN_25; 
  wire  _T_5_10; 
  wire  _GEN_26; 
  wire  _T_5_11; 
  wire  _GEN_27; 
  wire  _T_5_12; 
  wire  _GEN_28; 
  wire  _T_5_13; 
  wire  _GEN_29; 
  wire  _T_5_14; 
  wire  _GEN_30; 
  wire  _T_5_15; 
  wire  _GEN_31; 
  wire  _T_8; 
  wire  _T_10; 
  wire  _T_11; 
  wire [11:0] _T_6_0; 
  wire [11:0] _T_6_1; 
  wire [11:0] _GEN_33; 
  wire [11:0] _T_6_2; 
  wire [11:0] _GEN_34; 
  wire [11:0] _T_6_3; 
  wire [11:0] _GEN_35; 
  wire [11:0] _T_6_4; 
  wire [11:0] _GEN_36; 
  wire [11:0] _T_6_5; 
  wire [11:0] _GEN_37; 
  wire [11:0] _T_6_6; 
  wire [11:0] _GEN_38; 
  wire [11:0] _T_6_7; 
  wire [11:0] _GEN_39; 
  wire [11:0] _T_6_8; 
  wire [11:0] _GEN_40; 
  wire [11:0] _T_6_9; 
  wire [11:0] _GEN_41; 
  wire [11:0] _T_6_10; 
  wire [11:0] _GEN_42; 
  wire [11:0] _T_6_11; 
  wire [11:0] _GEN_43; 
  wire [11:0] _T_6_12; 
  wire [11:0] _GEN_44; 
  wire [11:0] _T_6_13; 
  wire [11:0] _GEN_45; 
  wire [11:0] _T_6_14; 
  wire [11:0] _GEN_46; 
  wire [11:0] _T_6_15; 
  wire [15:0] _T_13; 
  wire  _T_15; 
  wire  _T_16; 
  wire  _T_17; 
  wire  _T_18; 
  wire  _T_19; 
  wire  _T_20; 
  wire  _T_21; 
  wire  _T_22; 
  wire  _T_23; 
  wire  _T_24; 
  wire  _T_25; 
  wire  _T_26; 
  wire  _T_27; 
  wire  _T_28; 
  wire  _T_29; 
  wire  _T_30; 
  wire [15:0] _T_32; 
  wire  _T_34; 
  wire  _T_35; 
  wire  _T_36; 
  wire  _T_37; 
  wire  _T_38; 
  wire  _T_39; 
  wire  _T_40; 
  wire  _T_41; 
  wire  _T_42; 
  wire  _T_43; 
  wire  _T_44; 
  wire  _T_45; 
  wire  _T_46; 
  wire  _T_47; 
  wire  _T_48; 
  wire  _T_49; 
  wire  _T_50; 
  wire  _T_51; 
  wire  _T_53; 
  wire  _T_56; 
  wire  _T_61; 
  wire  _T_66; 
  wire  _T_71; 
  wire  _T_76; 
  wire  _T_81; 
  wire  _T_86; 
  wire  _T_91; 
  wire  _T_96; 
  wire  _T_101; 
  wire  _T_106; 
  wire  _T_111; 
  wire  _T_116; 
  wire  _T_121; 
  wire  _T_126; 
  wire  _T_130_0; 
  wire  _T_130_1; 
  wire  _GEN_49; 
  wire  _T_130_2; 
  wire  _GEN_50; 
  wire  _T_130_3; 
  wire  _GEN_51; 
  wire  _T_130_4; 
  wire  _GEN_52; 
  wire  _T_130_5; 
  wire  _GEN_53; 
  wire  _T_130_6; 
  wire  _GEN_54; 
  wire  _T_130_7; 
  wire  _GEN_55; 
  wire  _T_130_8; 
  wire  _GEN_56; 
  wire  _T_130_9; 
  wire  _GEN_57; 
  wire  _T_130_10; 
  wire  _GEN_58; 
  wire  _T_130_11; 
  wire  _GEN_59; 
  wire  _T_130_12; 
  wire  _GEN_60; 
  wire  _T_130_13; 
  wire  _GEN_61; 
  wire  _T_130_14; 
  wire  _GEN_62; 
  wire  _T_130_15; 
  wire  _GEN_63; 
  wire  _T_135; 
  wire  _T_133_0; 
  wire  _T_133_1; 
  wire  _GEN_65; 
  wire  _T_133_2; 
  wire  _GEN_66; 
  wire  _T_133_3; 
  wire  _GEN_67; 
  wire  _T_133_4; 
  wire  _GEN_68; 
  wire  _T_133_5; 
  wire  _GEN_69; 
  wire  _T_133_6; 
  wire  _GEN_70; 
  wire  _T_133_7; 
  wire  _GEN_71; 
  wire  _T_133_8; 
  wire  _GEN_72; 
  wire  _T_133_9; 
  wire  _GEN_73; 
  wire  _T_133_10; 
  wire  _GEN_74; 
  wire  _T_133_11; 
  wire  _GEN_75; 
  wire  _T_133_12; 
  wire  _GEN_76; 
  wire  _T_133_13; 
  wire  _GEN_77; 
  wire  _T_133_14; 
  wire  _GEN_78; 
  wire  _T_133_15; 
  wire  _GEN_79; 
  wire  _T_136; 
  wire  _T_138; 
  wire  _T_139; 
  wire [11:0] _T_134_0; 
  wire [11:0] _T_134_1; 
  wire [11:0] _GEN_81; 
  wire [11:0] _T_134_2; 
  wire [11:0] _GEN_82; 
  wire [11:0] _T_134_3; 
  wire [11:0] _GEN_83; 
  wire [11:0] _T_134_4; 
  wire [11:0] _GEN_84; 
  wire [11:0] _T_134_5; 
  wire [11:0] _GEN_85; 
  wire [11:0] _T_134_6; 
  wire [11:0] _GEN_86; 
  wire [11:0] _T_134_7; 
  wire [11:0] _GEN_87; 
  wire [11:0] _T_134_8; 
  wire [11:0] _GEN_88; 
  wire [11:0] _T_134_9; 
  wire [11:0] _GEN_89; 
  wire [11:0] _T_134_10; 
  wire [11:0] _GEN_90; 
  wire [11:0] _T_134_11; 
  wire [11:0] _GEN_91; 
  wire [11:0] _T_134_12; 
  wire [11:0] _GEN_92; 
  wire [11:0] _T_134_13; 
  wire [11:0] _GEN_93; 
  wire [11:0] _T_134_14; 
  wire [11:0] _GEN_94; 
  wire [11:0] _T_134_15; 
  wire [15:0] _T_141; 
  wire  _T_143; 
  wire  _T_144; 
  wire  _T_145; 
  wire  _T_146; 
  wire  _T_147; 
  wire  _T_148; 
  wire  _T_149; 
  wire  _T_150; 
  wire  _T_151; 
  wire  _T_152; 
  wire  _T_153; 
  wire  _T_154; 
  wire  _T_155; 
  wire  _T_156; 
  wire  _T_157; 
  wire  _T_158; 
  wire [15:0] _T_160; 
  wire  _T_162; 
  wire  _T_163; 
  wire  _T_164; 
  wire  _T_165; 
  wire  _T_166; 
  wire  _T_167; 
  wire  _T_168; 
  wire  _T_169; 
  wire  _T_170; 
  wire  _T_171; 
  wire  _T_172; 
  wire  _T_173; 
  wire  _T_174; 
  wire  _T_175; 
  wire  _T_176; 
  wire  _T_177; 
  wire  _T_178; 
  wire  _T_180; 
  dual_Queue_14 dual_Queue ( 
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits(Queue_io_enq_bits),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits(Queue_io_deq_bits)
  );
  dual_Queue_14 Queue_1 ( 
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits(Queue_1_io_enq_bits),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits(Queue_1_io_deq_bits)
  );
  dual_Queue_14 dual_Queue_2 ( 
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits(Queue_2_io_enq_bits),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits(Queue_2_io_deq_bits)
  );
  dual_Queue_14 Queue_3 ( 
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits(Queue_3_io_enq_bits),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits(Queue_3_io_deq_bits)
  );
  dual_Queue_14 dual_Queue_4 ( 
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits(Queue_4_io_enq_bits),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits(Queue_4_io_deq_bits)
  );
  dual_Queue_14 dual_Queue_5 ( 
    .clock(Queue_5_clock),
    .reset(Queue_5_reset),
    .io_enq_ready(Queue_5_io_enq_ready),
    .io_enq_valid(Queue_5_io_enq_valid),
    .io_enq_bits(Queue_5_io_enq_bits),
    .io_deq_ready(Queue_5_io_deq_ready),
    .io_deq_valid(Queue_5_io_deq_valid),
    .io_deq_bits(Queue_5_io_deq_bits)
  );
  dual_Queue_14 Queue_6 ( 
    .clock(Queue_6_clock),
    .reset(Queue_6_reset),
    .io_enq_ready(Queue_6_io_enq_ready),
    .io_enq_valid(Queue_6_io_enq_valid),
    .io_enq_bits(Queue_6_io_enq_bits),
    .io_deq_ready(Queue_6_io_deq_ready),
    .io_deq_valid(Queue_6_io_deq_valid),
    .io_deq_bits(Queue_6_io_deq_bits)
  );
  dual_Queue_21 Queue_7 ( 
    .clock(Queue_7_clock),
    .reset(Queue_7_reset),
    .io_enq_ready(Queue_7_io_enq_ready),
    .io_enq_valid(Queue_7_io_enq_valid),
    .io_enq_bits(Queue_7_io_enq_bits),
    .io_deq_ready(Queue_7_io_deq_ready),
    .io_deq_valid(Queue_7_io_deq_valid),
    .io_deq_bits(Queue_7_io_deq_bits)
  );
  dual_Queue_21 dual_Queue_8 ( 
    .clock(Queue_8_clock),
    .reset(Queue_8_reset),
    .io_enq_ready(Queue_8_io_enq_ready),
    .io_enq_valid(Queue_8_io_enq_valid),
    .io_enq_bits(Queue_8_io_enq_bits),
    .io_deq_ready(Queue_8_io_deq_ready),
    .io_deq_valid(Queue_8_io_deq_valid),
    .io_deq_bits(Queue_8_io_deq_bits)
  );
  dual_Queue_21 dual_Queue_9 ( 
    .clock(Queue_9_clock),
    .reset(Queue_9_reset),
    .io_enq_ready(Queue_9_io_enq_ready),
    .io_enq_valid(Queue_9_io_enq_valid),
    .io_enq_bits(Queue_9_io_enq_bits),
    .io_deq_ready(Queue_9_io_deq_ready),
    .io_deq_valid(Queue_9_io_deq_valid),
    .io_deq_bits(Queue_9_io_deq_bits)
  );
  dual_Queue_21 Queue_10 ( 
    .clock(Queue_10_clock),
    .reset(Queue_10_reset),
    .io_enq_ready(Queue_10_io_enq_ready),
    .io_enq_valid(Queue_10_io_enq_valid),
    .io_enq_bits(Queue_10_io_enq_bits),
    .io_deq_ready(Queue_10_io_deq_ready),
    .io_deq_valid(Queue_10_io_deq_valid),
    .io_deq_bits(Queue_10_io_deq_bits)
  );
  dual_Queue_21 Queue_11 ( 
    .clock(Queue_11_clock),
    .reset(Queue_11_reset),
    .io_enq_ready(Queue_11_io_enq_ready),
    .io_enq_valid(Queue_11_io_enq_valid),
    .io_enq_bits(Queue_11_io_enq_bits),
    .io_deq_ready(Queue_11_io_deq_ready),
    .io_deq_valid(Queue_11_io_deq_valid),
    .io_deq_bits(Queue_11_io_deq_bits)
  );
  dual_Queue_21 Queue_12 ( 
    .clock(Queue_12_clock),
    .reset(Queue_12_reset),
    .io_enq_ready(Queue_12_io_enq_ready),
    .io_enq_valid(Queue_12_io_enq_valid),
    .io_enq_bits(Queue_12_io_enq_bits),
    .io_deq_ready(Queue_12_io_deq_ready),
    .io_deq_valid(Queue_12_io_deq_valid),
    .io_deq_bits(Queue_12_io_deq_bits)
  );
  dual_Queue_21 Queue_13 ( 
    .clock(Queue_13_clock),
    .reset(Queue_13_reset),
    .io_enq_ready(Queue_13_io_enq_ready),
    .io_enq_valid(Queue_13_io_enq_valid),
    .io_enq_bits(Queue_13_io_enq_bits),
    .io_deq_ready(Queue_13_io_deq_ready),
    .io_deq_valid(Queue_13_io_deq_valid),
    .io_deq_bits(Queue_13_io_deq_bits)
  );
  dual_Queue_21 dual_Queue_14 ( 
    .clock(Queue_14_clock),
    .reset(Queue_14_reset),
    .io_enq_ready(Queue_14_io_enq_ready),
    .io_enq_valid(Queue_14_io_enq_valid),
    .io_enq_bits(Queue_14_io_enq_bits),
    .io_deq_ready(Queue_14_io_deq_ready),
    .io_deq_valid(Queue_14_io_deq_valid),
    .io_deq_bits(Queue_14_io_deq_bits)
  );
  dual_Queue_21 Queue_15 ( 
    .clock(Queue_15_clock),
    .reset(Queue_15_reset),
    .io_enq_ready(Queue_15_io_enq_ready),
    .io_enq_valid(Queue_15_io_enq_valid),
    .io_enq_bits(Queue_15_io_enq_bits),
    .io_deq_ready(Queue_15_io_deq_ready),
    .io_deq_valid(Queue_15_io_deq_valid),
    .io_deq_bits(Queue_15_io_deq_bits)
  );
  dual_Queue_14 Queue_16 ( 
    .clock(Queue_16_clock),
    .reset(Queue_16_reset),
    .io_enq_ready(Queue_16_io_enq_ready),
    .io_enq_valid(Queue_16_io_enq_valid),
    .io_enq_bits(Queue_16_io_enq_bits),
    .io_deq_ready(Queue_16_io_deq_ready),
    .io_deq_valid(Queue_16_io_deq_valid),
    .io_deq_bits(Queue_16_io_deq_bits)
  );
  dual_Queue_14 Queue_17 ( 
    .clock(Queue_17_clock),
    .reset(Queue_17_reset),
    .io_enq_ready(Queue_17_io_enq_ready),
    .io_enq_valid(Queue_17_io_enq_valid),
    .io_enq_bits(Queue_17_io_enq_bits),
    .io_deq_ready(Queue_17_io_deq_ready),
    .io_deq_valid(Queue_17_io_deq_valid),
    .io_deq_bits(Queue_17_io_deq_bits)
  );
  dual_Queue_14 Queue_18 ( 
    .clock(Queue_18_clock),
    .reset(Queue_18_reset),
    .io_enq_ready(Queue_18_io_enq_ready),
    .io_enq_valid(Queue_18_io_enq_valid),
    .io_enq_bits(Queue_18_io_enq_bits),
    .io_deq_ready(Queue_18_io_deq_ready),
    .io_deq_valid(Queue_18_io_deq_valid),
    .io_deq_bits(Queue_18_io_deq_bits)
  );
  dual_Queue_14 Queue_19 ( 
    .clock(Queue_19_clock),
    .reset(Queue_19_reset),
    .io_enq_ready(Queue_19_io_enq_ready),
    .io_enq_valid(Queue_19_io_enq_valid),
    .io_enq_bits(Queue_19_io_enq_bits),
    .io_deq_ready(Queue_19_io_deq_ready),
    .io_deq_valid(Queue_19_io_deq_valid),
    .io_deq_bits(Queue_19_io_deq_bits)
  );
  dual_Queue_14 Queue_20 ( 
    .clock(Queue_20_clock),
    .reset(Queue_20_reset),
    .io_enq_ready(Queue_20_io_enq_ready),
    .io_enq_valid(Queue_20_io_enq_valid),
    .io_enq_bits(Queue_20_io_enq_bits),
    .io_deq_ready(Queue_20_io_deq_ready),
    .io_deq_valid(Queue_20_io_deq_valid),
    .io_deq_bits(Queue_20_io_deq_bits)
  );
  dual_Queue_14 dual_Queue_21 ( 
    .clock(Queue_21_clock),
    .reset(Queue_21_reset),
    .io_enq_ready(Queue_21_io_enq_ready),
    .io_enq_valid(Queue_21_io_enq_valid),
    .io_enq_bits(Queue_21_io_enq_bits),
    .io_deq_ready(Queue_21_io_deq_ready),
    .io_deq_valid(Queue_21_io_deq_valid),
    .io_deq_bits(Queue_21_io_deq_bits)
  );
  dual_Queue_14 Queue_22 ( 
    .clock(Queue_22_clock),
    .reset(Queue_22_reset),
    .io_enq_ready(Queue_22_io_enq_ready),
    .io_enq_valid(Queue_22_io_enq_valid),
    .io_enq_bits(Queue_22_io_enq_bits),
    .io_deq_ready(Queue_22_io_deq_ready),
    .io_deq_valid(Queue_22_io_deq_valid),
    .io_deq_bits(Queue_22_io_deq_bits)
  );
  dual_Queue_21 Queue_23 ( 
    .clock(Queue_23_clock),
    .reset(Queue_23_reset),
    .io_enq_ready(Queue_23_io_enq_ready),
    .io_enq_valid(Queue_23_io_enq_valid),
    .io_enq_bits(Queue_23_io_enq_bits),
    .io_deq_ready(Queue_23_io_deq_ready),
    .io_deq_valid(Queue_23_io_deq_valid),
    .io_deq_bits(Queue_23_io_deq_bits)
  );
  dual_Queue_21 Queue_24 ( 
    .clock(Queue_24_clock),
    .reset(Queue_24_reset),
    .io_enq_ready(Queue_24_io_enq_ready),
    .io_enq_valid(Queue_24_io_enq_valid),
    .io_enq_bits(Queue_24_io_enq_bits),
    .io_deq_ready(Queue_24_io_deq_ready),
    .io_deq_valid(Queue_24_io_deq_valid),
    .io_deq_bits(Queue_24_io_deq_bits)
  );
  dual_Queue_21 Queue_25 ( 
    .clock(Queue_25_clock),
    .reset(Queue_25_reset),
    .io_enq_ready(Queue_25_io_enq_ready),
    .io_enq_valid(Queue_25_io_enq_valid),
    .io_enq_bits(Queue_25_io_enq_bits),
    .io_deq_ready(Queue_25_io_deq_ready),
    .io_deq_valid(Queue_25_io_deq_valid),
    .io_deq_bits(Queue_25_io_deq_bits)
  );
  dual_Queue_21 Queue_26 ( 
    .clock(Queue_26_clock),
    .reset(Queue_26_reset),
    .io_enq_ready(Queue_26_io_enq_ready),
    .io_enq_valid(Queue_26_io_enq_valid),
    .io_enq_bits(Queue_26_io_enq_bits),
    .io_deq_ready(Queue_26_io_deq_ready),
    .io_deq_valid(Queue_26_io_deq_valid),
    .io_deq_bits(Queue_26_io_deq_bits)
  );
  dual_Queue_21 Queue_27 ( 
    .clock(Queue_27_clock),
    .reset(Queue_27_reset),
    .io_enq_ready(Queue_27_io_enq_ready),
    .io_enq_valid(Queue_27_io_enq_valid),
    .io_enq_bits(Queue_27_io_enq_bits),
    .io_deq_ready(Queue_27_io_deq_ready),
    .io_deq_valid(Queue_27_io_deq_valid),
    .io_deq_bits(Queue_27_io_deq_bits)
  );
  dual_Queue_21 Queue_28 ( 
    .clock(Queue_28_clock),
    .reset(Queue_28_reset),
    .io_enq_ready(Queue_28_io_enq_ready),
    .io_enq_valid(Queue_28_io_enq_valid),
    .io_enq_bits(Queue_28_io_enq_bits),
    .io_deq_ready(Queue_28_io_deq_ready),
    .io_deq_valid(Queue_28_io_deq_valid),
    .io_deq_bits(Queue_28_io_deq_bits)
  );
  dual_Queue_21 Queue_29 ( 
    .clock(Queue_29_clock),
    .reset(Queue_29_reset),
    .io_enq_ready(Queue_29_io_enq_ready),
    .io_enq_valid(Queue_29_io_enq_valid),
    .io_enq_bits(Queue_29_io_enq_bits),
    .io_deq_ready(Queue_29_io_deq_ready),
    .io_deq_valid(Queue_29_io_deq_valid),
    .io_deq_bits(Queue_29_io_deq_bits)
  );
  dual_Queue_21 Queue_30 ( 
    .clock(Queue_30_clock),
    .reset(Queue_30_reset),
    .io_enq_ready(Queue_30_io_enq_ready),
    .io_enq_valid(Queue_30_io_enq_valid),
    .io_enq_bits(Queue_30_io_enq_bits),
    .io_deq_ready(Queue_30_io_deq_ready),
    .io_deq_valid(Queue_30_io_deq_valid),
    .io_deq_bits(Queue_30_io_deq_bits)
  );
  dual_Queue_21 Queue_31 ( 
    .clock(Queue_31_clock),
    .reset(Queue_31_reset),
    .io_enq_ready(Queue_31_io_enq_ready),
    .io_enq_valid(Queue_31_io_enq_valid),
    .io_enq_bits(Queue_31_io_enq_bits),
    .io_deq_ready(Queue_31_io_deq_ready),
    .io_deq_valid(Queue_31_io_deq_valid),
    .io_deq_bits(Queue_31_io_deq_bits)
  );
  assign _T_2_0 = Queue_io_enq_ready; 
  assign _T_2_1 = Queue_1_io_enq_ready; 
  assign _GEN_1 = 4'h1 == auto_in_arid ? _T_2_1 : _T_2_0; 
  assign _T_2_2 = Queue_2_io_enq_ready; 
  assign _GEN_2 = 4'h2 == auto_in_arid ? _T_2_2 : _GEN_1; 
  assign _T_2_3 = Queue_3_io_enq_ready; 
  assign _GEN_3 = 4'h3 == auto_in_arid ? _T_2_3 : _GEN_2; 
  assign _T_2_4 = Queue_4_io_enq_ready; 
  assign _GEN_4 = 4'h4 == auto_in_arid ? _T_2_4 : _GEN_3; 
  assign _T_2_5 = Queue_5_io_enq_ready; 
  assign _GEN_5 = 4'h5 == auto_in_arid ? _T_2_5 : _GEN_4; 
  assign _T_2_6 = Queue_6_io_enq_ready; 
  assign _GEN_6 = 4'h6 == auto_in_arid ? _T_2_6 : _GEN_5; 
  assign _T_2_7 = Queue_7_io_enq_ready; 
  assign _GEN_7 = 4'h7 == auto_in_arid ? _T_2_7 : _GEN_6; 
  assign _T_2_8 = Queue_8_io_enq_ready; 
  assign _GEN_8 = 4'h8 == auto_in_arid ? _T_2_8 : _GEN_7; 
  assign _T_2_9 = Queue_9_io_enq_ready; 
  assign _GEN_9 = 4'h9 == auto_in_arid ? _T_2_9 : _GEN_8; 
  assign _T_2_10 = Queue_10_io_enq_ready; 
  assign _GEN_10 = 4'ha == auto_in_arid ? _T_2_10 : _GEN_9; 
  assign _T_2_11 = Queue_11_io_enq_ready; 
  assign _GEN_11 = 4'hb == auto_in_arid ? _T_2_11 : _GEN_10; 
  assign _T_2_12 = Queue_12_io_enq_ready; 
  assign _GEN_12 = 4'hc == auto_in_arid ? _T_2_12 : _GEN_11; 
  assign _T_2_13 = Queue_13_io_enq_ready; 
  assign _GEN_13 = 4'hd == auto_in_arid ? _T_2_13 : _GEN_12; 
  assign _T_2_14 = Queue_14_io_enq_ready; 
  assign _GEN_14 = 4'he == auto_in_arid ? _T_2_14 : _GEN_13; 
  assign _T_2_15 = Queue_15_io_enq_ready; 
  assign _GEN_15 = 4'hf == auto_in_arid ? _T_2_15 : _GEN_14; 
  assign _T_7 = auto_out_rvalid == 1'h0; 
  assign _T_5_0 = Queue_io_deq_valid; 
  assign _T_5_1 = Queue_1_io_deq_valid; 
  assign _GEN_17 = 4'h1 == auto_out_rid ? _T_5_1 : _T_5_0; 
  assign _T_5_2 = Queue_2_io_deq_valid; 
  assign _GEN_18 = 4'h2 == auto_out_rid ? _T_5_2 : _GEN_17; 
  assign _T_5_3 = Queue_3_io_deq_valid; 
  assign _GEN_19 = 4'h3 == auto_out_rid ? _T_5_3 : _GEN_18; 
  assign _T_5_4 = Queue_4_io_deq_valid; 
  assign _GEN_20 = 4'h4 == auto_out_rid ? _T_5_4 : _GEN_19; 
  assign _T_5_5 = Queue_5_io_deq_valid; 
  assign _GEN_21 = 4'h5 == auto_out_rid ? _T_5_5 : _GEN_20; 
  assign _T_5_6 = Queue_6_io_deq_valid; 
  assign _GEN_22 = 4'h6 == auto_out_rid ? _T_5_6 : _GEN_21; 
  assign _T_5_7 = Queue_7_io_deq_valid; 
  assign _GEN_23 = 4'h7 == auto_out_rid ? _T_5_7 : _GEN_22; 
  assign _T_5_8 = Queue_8_io_deq_valid; 
  assign _GEN_24 = 4'h8 == auto_out_rid ? _T_5_8 : _GEN_23; 
  assign _T_5_9 = Queue_9_io_deq_valid; 
  assign _GEN_25 = 4'h9 == auto_out_rid ? _T_5_9 : _GEN_24; 
  assign _T_5_10 = Queue_10_io_deq_valid; 
  assign _GEN_26 = 4'ha == auto_out_rid ? _T_5_10 : _GEN_25; 
  assign _T_5_11 = Queue_11_io_deq_valid; 
  assign _GEN_27 = 4'hb == auto_out_rid ? _T_5_11 : _GEN_26; 
  assign _T_5_12 = Queue_12_io_deq_valid; 
  assign _GEN_28 = 4'hc == auto_out_rid ? _T_5_12 : _GEN_27; 
  assign _T_5_13 = Queue_13_io_deq_valid; 
  assign _GEN_29 = 4'hd == auto_out_rid ? _T_5_13 : _GEN_28; 
  assign _T_5_14 = Queue_14_io_deq_valid; 
  assign _GEN_30 = 4'he == auto_out_rid ? _T_5_14 : _GEN_29; 
  assign _T_5_15 = Queue_15_io_deq_valid; 
  assign _GEN_31 = 4'hf == auto_out_rid ? _T_5_15 : _GEN_30; 
  assign _T_8 = _T_7 | _GEN_31; 
  assign _T_10 = _T_8 | reset; 
  assign _T_11 = _T_10 == 1'h0; 
  assign _T_6_0 = Queue_io_deq_bits; 
  assign _T_6_1 = Queue_1_io_deq_bits; 
  assign _GEN_33 = 4'h1 == auto_out_rid ? _T_6_1 : _T_6_0; 
  assign _T_6_2 = Queue_2_io_deq_bits; 
  assign _GEN_34 = 4'h2 == auto_out_rid ? _T_6_2 : _GEN_33; 
  assign _T_6_3 = Queue_3_io_deq_bits; 
  assign _GEN_35 = 4'h3 == auto_out_rid ? _T_6_3 : _GEN_34; 
  assign _T_6_4 = Queue_4_io_deq_bits; 
  assign _GEN_36 = 4'h4 == auto_out_rid ? _T_6_4 : _GEN_35; 
  assign _T_6_5 = Queue_5_io_deq_bits; 
  assign _GEN_37 = 4'h5 == auto_out_rid ? _T_6_5 : _GEN_36; 
  assign _T_6_6 = Queue_6_io_deq_bits; 
  assign _GEN_38 = 4'h6 == auto_out_rid ? _T_6_6 : _GEN_37; 
  assign _T_6_7 = Queue_7_io_deq_bits; 
  assign _GEN_39 = 4'h7 == auto_out_rid ? _T_6_7 : _GEN_38; 
  assign _T_6_8 = Queue_8_io_deq_bits; 
  assign _GEN_40 = 4'h8 == auto_out_rid ? _T_6_8 : _GEN_39; 
  assign _T_6_9 = Queue_9_io_deq_bits; 
  assign _GEN_41 = 4'h9 == auto_out_rid ? _T_6_9 : _GEN_40; 
  assign _T_6_10 = Queue_10_io_deq_bits; 
  assign _GEN_42 = 4'ha == auto_out_rid ? _T_6_10 : _GEN_41; 
  assign _T_6_11 = Queue_11_io_deq_bits; 
  assign _GEN_43 = 4'hb == auto_out_rid ? _T_6_11 : _GEN_42; 
  assign _T_6_12 = Queue_12_io_deq_bits; 
  assign _GEN_44 = 4'hc == auto_out_rid ? _T_6_12 : _GEN_43; 
  assign _T_6_13 = Queue_13_io_deq_bits; 
  assign _GEN_45 = 4'hd == auto_out_rid ? _T_6_13 : _GEN_44; 
  assign _T_6_14 = Queue_14_io_deq_bits; 
  assign _GEN_46 = 4'he == auto_out_rid ? _T_6_14 : _GEN_45; 
  assign _T_6_15 = Queue_15_io_deq_bits; 
  assign _T_13 = 16'h1 << auto_in_arid; 
  assign _T_15 = _T_13[0]; 
  assign _T_16 = _T_13[1]; 
  assign _T_17 = _T_13[2]; 
  assign _T_18 = _T_13[3]; 
  assign _T_19 = _T_13[4]; 
  assign _T_20 = _T_13[5]; 
  assign _T_21 = _T_13[6]; 
  assign _T_22 = _T_13[7]; 
  assign _T_23 = _T_13[8]; 
  assign _T_24 = _T_13[9]; 
  assign _T_25 = _T_13[10]; 
  assign _T_26 = _T_13[11]; 
  assign _T_27 = _T_13[12]; 
  assign _T_28 = _T_13[13]; 
  assign _T_29 = _T_13[14]; 
  assign _T_30 = _T_13[15]; 
  assign _T_32 = 16'h1 << auto_out_rid; 
  assign _T_34 = _T_32[0]; 
  assign _T_35 = _T_32[1]; 
  assign _T_36 = _T_32[2]; 
  assign _T_37 = _T_32[3]; 
  assign _T_38 = _T_32[4]; 
  assign _T_39 = _T_32[5]; 
  assign _T_40 = _T_32[6]; 
  assign _T_41 = _T_32[7]; 
  assign _T_42 = _T_32[8]; 
  assign _T_43 = _T_32[9]; 
  assign _T_44 = _T_32[10]; 
  assign _T_45 = _T_32[11]; 
  assign _T_46 = _T_32[12]; 
  assign _T_47 = _T_32[13]; 
  assign _T_48 = _T_32[14]; 
  assign _T_49 = _T_32[15]; 
  assign _T_50 = auto_out_rvalid & auto_in_rready; 
  assign _T_51 = _T_50 & _T_34; 
  assign _T_53 = auto_in_arvalid & auto_out_arready; 
  assign _T_56 = _T_50 & _T_35; 
  assign _T_61 = _T_50 & _T_36; 
  assign _T_66 = _T_50 & _T_37; 
  assign _T_71 = _T_50 & _T_38; 
  assign _T_76 = _T_50 & _T_39; 
  assign _T_81 = _T_50 & _T_40; 
  assign _T_86 = _T_50 & _T_41; 
  assign _T_91 = _T_50 & _T_42; 
  assign _T_96 = _T_50 & _T_43; 
  assign _T_101 = _T_50 & _T_44; 
  assign _T_106 = _T_50 & _T_45; 
  assign _T_111 = _T_50 & _T_46; 
  assign _T_116 = _T_50 & _T_47; 
  assign _T_121 = _T_50 & _T_48; 
  assign _T_126 = _T_50 & _T_49; 
  assign _T_130_0 = Queue_16_io_enq_ready; 
  assign _T_130_1 = Queue_17_io_enq_ready; 
  assign _GEN_49 = 4'h1 == auto_in_awid ? _T_130_1 : _T_130_0; 
  assign _T_130_2 = Queue_18_io_enq_ready; 
  assign _GEN_50 = 4'h2 == auto_in_awid ? _T_130_2 : _GEN_49; 
  assign _T_130_3 = Queue_19_io_enq_ready; 
  assign _GEN_51 = 4'h3 == auto_in_awid ? _T_130_3 : _GEN_50; 
  assign _T_130_4 = Queue_20_io_enq_ready; 
  assign _GEN_52 = 4'h4 == auto_in_awid ? _T_130_4 : _GEN_51; 
  assign _T_130_5 = Queue_21_io_enq_ready; 
  assign _GEN_53 = 4'h5 == auto_in_awid ? _T_130_5 : _GEN_52; 
  assign _T_130_6 = Queue_22_io_enq_ready; 
  assign _GEN_54 = 4'h6 == auto_in_awid ? _T_130_6 : _GEN_53; 
  assign _T_130_7 = Queue_23_io_enq_ready; 
  assign _GEN_55 = 4'h7 == auto_in_awid ? _T_130_7 : _GEN_54; 
  assign _T_130_8 = Queue_24_io_enq_ready; 
  assign _GEN_56 = 4'h8 == auto_in_awid ? _T_130_8 : _GEN_55; 
  assign _T_130_9 = Queue_25_io_enq_ready; 
  assign _GEN_57 = 4'h9 == auto_in_awid ? _T_130_9 : _GEN_56; 
  assign _T_130_10 = Queue_26_io_enq_ready; 
  assign _GEN_58 = 4'ha == auto_in_awid ? _T_130_10 : _GEN_57; 
  assign _T_130_11 = Queue_27_io_enq_ready; 
  assign _GEN_59 = 4'hb == auto_in_awid ? _T_130_11 : _GEN_58; 
  assign _T_130_12 = Queue_28_io_enq_ready; 
  assign _GEN_60 = 4'hc == auto_in_awid ? _T_130_12 : _GEN_59; 
  assign _T_130_13 = Queue_29_io_enq_ready; 
  assign _GEN_61 = 4'hd == auto_in_awid ? _T_130_13 : _GEN_60; 
  assign _T_130_14 = Queue_30_io_enq_ready; 
  assign _GEN_62 = 4'he == auto_in_awid ? _T_130_14 : _GEN_61; 
  assign _T_130_15 = Queue_31_io_enq_ready; 
  assign _GEN_63 = 4'hf == auto_in_awid ? _T_130_15 : _GEN_62; 
  assign _T_135 = auto_out_bvalid == 1'h0; 
  assign _T_133_0 = Queue_16_io_deq_valid; 
  assign _T_133_1 = Queue_17_io_deq_valid; 
  assign _GEN_65 = 4'h1 == auto_out_bid ? _T_133_1 : _T_133_0; 
  assign _T_133_2 = Queue_18_io_deq_valid; 
  assign _GEN_66 = 4'h2 == auto_out_bid ? _T_133_2 : _GEN_65; 
  assign _T_133_3 = Queue_19_io_deq_valid; 
  assign _GEN_67 = 4'h3 == auto_out_bid ? _T_133_3 : _GEN_66; 
  assign _T_133_4 = Queue_20_io_deq_valid; 
  assign _GEN_68 = 4'h4 == auto_out_bid ? _T_133_4 : _GEN_67; 
  assign _T_133_5 = Queue_21_io_deq_valid; 
  assign _GEN_69 = 4'h5 == auto_out_bid ? _T_133_5 : _GEN_68; 
  assign _T_133_6 = Queue_22_io_deq_valid; 
  assign _GEN_70 = 4'h6 == auto_out_bid ? _T_133_6 : _GEN_69; 
  assign _T_133_7 = Queue_23_io_deq_valid; 
  assign _GEN_71 = 4'h7 == auto_out_bid ? _T_133_7 : _GEN_70; 
  assign _T_133_8 = Queue_24_io_deq_valid; 
  assign _GEN_72 = 4'h8 == auto_out_bid ? _T_133_8 : _GEN_71; 
  assign _T_133_9 = Queue_25_io_deq_valid; 
  assign _GEN_73 = 4'h9 == auto_out_bid ? _T_133_9 : _GEN_72; 
  assign _T_133_10 = Queue_26_io_deq_valid; 
  assign _GEN_74 = 4'ha == auto_out_bid ? _T_133_10 : _GEN_73; 
  assign _T_133_11 = Queue_27_io_deq_valid; 
  assign _GEN_75 = 4'hb == auto_out_bid ? _T_133_11 : _GEN_74; 
  assign _T_133_12 = Queue_28_io_deq_valid; 
  assign _GEN_76 = 4'hc == auto_out_bid ? _T_133_12 : _GEN_75; 
  assign _T_133_13 = Queue_29_io_deq_valid; 
  assign _GEN_77 = 4'hd == auto_out_bid ? _T_133_13 : _GEN_76; 
  assign _T_133_14 = Queue_30_io_deq_valid; 
  assign _GEN_78 = 4'he == auto_out_bid ? _T_133_14 : _GEN_77; 
  assign _T_133_15 = Queue_31_io_deq_valid; 
  assign _GEN_79 = 4'hf == auto_out_bid ? _T_133_15 : _GEN_78; 
  assign _T_136 = _T_135 | _GEN_79; 
  assign _T_138 = _T_136 | reset; 
  assign _T_139 = _T_138 == 1'h0; 
  assign _T_134_0 = Queue_16_io_deq_bits; 
  assign _T_134_1 = Queue_17_io_deq_bits; 
  assign _GEN_81 = 4'h1 == auto_out_bid ? _T_134_1 : _T_134_0; 
  assign _T_134_2 = Queue_18_io_deq_bits; 
  assign _GEN_82 = 4'h2 == auto_out_bid ? _T_134_2 : _GEN_81; 
  assign _T_134_3 = Queue_19_io_deq_bits; 
  assign _GEN_83 = 4'h3 == auto_out_bid ? _T_134_3 : _GEN_82; 
  assign _T_134_4 = Queue_20_io_deq_bits; 
  assign _GEN_84 = 4'h4 == auto_out_bid ? _T_134_4 : _GEN_83; 
  assign _T_134_5 = Queue_21_io_deq_bits; 
  assign _GEN_85 = 4'h5 == auto_out_bid ? _T_134_5 : _GEN_84; 
  assign _T_134_6 = Queue_22_io_deq_bits; 
  assign _GEN_86 = 4'h6 == auto_out_bid ? _T_134_6 : _GEN_85; 
  assign _T_134_7 = Queue_23_io_deq_bits; 
  assign _GEN_87 = 4'h7 == auto_out_bid ? _T_134_7 : _GEN_86; 
  assign _T_134_8 = Queue_24_io_deq_bits; 
  assign _GEN_88 = 4'h8 == auto_out_bid ? _T_134_8 : _GEN_87; 
  assign _T_134_9 = Queue_25_io_deq_bits; 
  assign _GEN_89 = 4'h9 == auto_out_bid ? _T_134_9 : _GEN_88; 
  assign _T_134_10 = Queue_26_io_deq_bits; 
  assign _GEN_90 = 4'ha == auto_out_bid ? _T_134_10 : _GEN_89; 
  assign _T_134_11 = Queue_27_io_deq_bits; 
  assign _GEN_91 = 4'hb == auto_out_bid ? _T_134_11 : _GEN_90; 
  assign _T_134_12 = Queue_28_io_deq_bits; 
  assign _GEN_92 = 4'hc == auto_out_bid ? _T_134_12 : _GEN_91; 
  assign _T_134_13 = Queue_29_io_deq_bits; 
  assign _GEN_93 = 4'hd == auto_out_bid ? _T_134_13 : _GEN_92; 
  assign _T_134_14 = Queue_30_io_deq_bits; 
  assign _GEN_94 = 4'he == auto_out_bid ? _T_134_14 : _GEN_93; 
  assign _T_134_15 = Queue_31_io_deq_bits; 
  assign _T_141 = 16'h1 << auto_in_awid; 
  assign _T_143 = _T_141[0]; 
  assign _T_144 = _T_141[1]; 
  assign _T_145 = _T_141[2]; 
  assign _T_146 = _T_141[3]; 
  assign _T_147 = _T_141[4]; 
  assign _T_148 = _T_141[5]; 
  assign _T_149 = _T_141[6]; 
  assign _T_150 = _T_141[7]; 
  assign _T_151 = _T_141[8]; 
  assign _T_152 = _T_141[9]; 
  assign _T_153 = _T_141[10]; 
  assign _T_154 = _T_141[11]; 
  assign _T_155 = _T_141[12]; 
  assign _T_156 = _T_141[13]; 
  assign _T_157 = _T_141[14]; 
  assign _T_158 = _T_141[15]; 
  assign _T_160 = 16'h1 << auto_out_bid; 
  assign _T_162 = _T_160[0]; 
  assign _T_163 = _T_160[1]; 
  assign _T_164 = _T_160[2]; 
  assign _T_165 = _T_160[3]; 
  assign _T_166 = _T_160[4]; 
  assign _T_167 = _T_160[5]; 
  assign _T_168 = _T_160[6]; 
  assign _T_169 = _T_160[7]; 
  assign _T_170 = _T_160[8]; 
  assign _T_171 = _T_160[9]; 
  assign _T_172 = _T_160[10]; 
  assign _T_173 = _T_160[11]; 
  assign _T_174 = _T_160[12]; 
  assign _T_175 = _T_160[13]; 
  assign _T_176 = _T_160[14]; 
  assign _T_177 = _T_160[15]; 
  assign _T_178 = auto_out_bvalid & auto_in_bready; 
  assign _T_180 = auto_in_awvalid & auto_out_awready; 
  assign auto_in_awready = auto_out_awready & _GEN_63; 
  assign auto_in_wready = auto_out_wready; 
  assign auto_in_bvalid = auto_out_bvalid; 
  assign auto_in_bid = auto_out_bid; 
  assign auto_in_bresp = auto_out_bresp; 
  assign auto_in_buser = 4'hf == auto_out_bid ? _T_134_15 : _GEN_94; 
  assign auto_in_arready = auto_out_arready & _GEN_15; 
  assign auto_in_rvalid = auto_out_rvalid; 
  assign auto_in_rid = auto_out_rid; 
  assign auto_in_rdata = auto_out_rdata; 
  assign auto_in_rresp = auto_out_rresp; 
  assign auto_in_ruser = 4'hf == auto_out_rid ? _T_6_15 : _GEN_46; 
  assign auto_in_rlast = auto_out_rlast; 
  assign auto_out_awvalid = auto_in_awvalid & _GEN_63; 
  assign auto_out_awid = auto_in_awid; 
  assign auto_out_awaddr = auto_in_awaddr; 
  assign auto_out_awlen = auto_in_awlen; 
  assign auto_out_awsize = auto_in_awsize; 
  assign auto_out_awburst = auto_in_awburst; 
  assign auto_out_awlock = auto_in_awlock; 
  assign auto_out_awcache = auto_in_awcache; 
  assign auto_out_awprot = auto_in_awprot; 
  assign auto_out_awqos = auto_in_awqos; 
  assign auto_out_awinstret = auto_in_awinstret; 
  assign auto_out_wvalid = auto_in_wvalid; 
  assign auto_out_wdata = auto_in_wdata; 
  assign auto_out_wstrb = auto_in_wstrb; 
  assign auto_out_wlast = auto_in_wlast; 
  assign auto_out_bready = auto_in_bready; 
  assign auto_out_arvalid = auto_in_arvalid & _GEN_15; 
  assign auto_out_arid = auto_in_arid; 
  assign auto_out_araddr = auto_in_araddr; 
  assign auto_out_arlen = auto_in_arlen; 
  assign auto_out_arsize = auto_in_arsize; 
  assign auto_out_arburst = auto_in_arburst; 
  assign auto_out_arlock = auto_in_arlock; 
  assign auto_out_arcache = auto_in_arcache; 
  assign auto_out_arprot = auto_in_arprot; 
  assign auto_out_arqos = auto_in_arqos; 
  assign auto_out_arinstret = auto_in_arinstret; 
  assign auto_out_rready = auto_in_rready; 
  assign Queue_clock = clock; 
  assign Queue_reset = reset; 
  assign Queue_io_enq_valid = _T_53 & _T_15; 
  assign Queue_io_enq_bits = auto_in_aruser; 
  assign Queue_io_deq_ready = _T_51 & auto_out_rlast; 
  assign Queue_1_clock = clock; 
  assign Queue_1_reset = reset; 
  assign Queue_1_io_enq_valid = _T_53 & _T_16; 
  assign Queue_1_io_enq_bits = auto_in_aruser; 
  assign Queue_1_io_deq_ready = _T_56 & auto_out_rlast; 
  assign Queue_2_clock = clock; 
  assign Queue_2_reset = reset; 
  assign Queue_2_io_enq_valid = _T_53 & _T_17; 
  assign Queue_2_io_enq_bits = auto_in_aruser; 
  assign Queue_2_io_deq_ready = _T_61 & auto_out_rlast; 
  assign Queue_3_clock = clock; 
  assign Queue_3_reset = reset; 
  assign Queue_3_io_enq_valid = _T_53 & _T_18; 
  assign Queue_3_io_enq_bits = auto_in_aruser; 
  assign Queue_3_io_deq_ready = _T_66 & auto_out_rlast; 
  assign Queue_4_clock = clock; 
  assign Queue_4_reset = reset; 
  assign Queue_4_io_enq_valid = _T_53 & _T_19; 
  assign Queue_4_io_enq_bits = auto_in_aruser; 
  assign Queue_4_io_deq_ready = _T_71 & auto_out_rlast; 
  assign Queue_5_clock = clock; 
  assign Queue_5_reset = reset; 
  assign Queue_5_io_enq_valid = _T_53 & _T_20; 
  assign Queue_5_io_enq_bits = auto_in_aruser; 
  assign Queue_5_io_deq_ready = _T_76 & auto_out_rlast; 
  assign Queue_6_clock = clock; 
  assign Queue_6_reset = reset; 
  assign Queue_6_io_enq_valid = _T_53 & _T_21; 
  assign Queue_6_io_enq_bits = auto_in_aruser; 
  assign Queue_6_io_deq_ready = _T_81 & auto_out_rlast; 
  assign Queue_7_clock = clock; 
  assign Queue_7_reset = reset; 
  assign Queue_7_io_enq_valid = _T_53 & _T_22; 
  assign Queue_7_io_enq_bits = auto_in_aruser; 
  assign Queue_7_io_deq_ready = _T_86 & auto_out_rlast; 
  assign Queue_8_clock = clock; 
  assign Queue_8_reset = reset; 
  assign Queue_8_io_enq_valid = _T_53 & _T_23; 
  assign Queue_8_io_enq_bits = auto_in_aruser; 
  assign Queue_8_io_deq_ready = _T_91 & auto_out_rlast; 
  assign Queue_9_clock = clock; 
  assign Queue_9_reset = reset; 
  assign Queue_9_io_enq_valid = _T_53 & _T_24; 
  assign Queue_9_io_enq_bits = auto_in_aruser; 
  assign Queue_9_io_deq_ready = _T_96 & auto_out_rlast; 
  assign Queue_10_clock = clock; 
  assign Queue_10_reset = reset; 
  assign Queue_10_io_enq_valid = _T_53 & _T_25; 
  assign Queue_10_io_enq_bits = auto_in_aruser; 
  assign Queue_10_io_deq_ready = _T_101 & auto_out_rlast; 
  assign Queue_11_clock = clock; 
  assign Queue_11_reset = reset; 
  assign Queue_11_io_enq_valid = _T_53 & _T_26; 
  assign Queue_11_io_enq_bits = auto_in_aruser; 
  assign Queue_11_io_deq_ready = _T_106 & auto_out_rlast; 
  assign Queue_12_clock = clock; 
  assign Queue_12_reset = reset; 
  assign Queue_12_io_enq_valid = _T_53 & _T_27; 
  assign Queue_12_io_enq_bits = auto_in_aruser; 
  assign Queue_12_io_deq_ready = _T_111 & auto_out_rlast; 
  assign Queue_13_clock = clock; 
  assign Queue_13_reset = reset; 
  assign Queue_13_io_enq_valid = _T_53 & _T_28; 
  assign Queue_13_io_enq_bits = auto_in_aruser; 
  assign Queue_13_io_deq_ready = _T_116 & auto_out_rlast; 
  assign Queue_14_clock = clock; 
  assign Queue_14_reset = reset; 
  assign Queue_14_io_enq_valid = _T_53 & _T_29; 
  assign Queue_14_io_enq_bits = auto_in_aruser; 
  assign Queue_14_io_deq_ready = _T_121 & auto_out_rlast; 
  assign Queue_15_clock = clock; 
  assign Queue_15_reset = reset; 
  assign Queue_15_io_enq_valid = _T_53 & _T_30; 
  assign Queue_15_io_enq_bits = auto_in_aruser; 
  assign Queue_15_io_deq_ready = _T_126 & auto_out_rlast; 
  assign Queue_16_clock = clock; 
  assign Queue_16_reset = reset; 
  assign Queue_16_io_enq_valid = _T_180 & _T_143; 
  assign Queue_16_io_enq_bits = auto_in_awuser; 
  assign Queue_16_io_deq_ready = _T_178 & _T_162; 
  assign Queue_17_clock = clock; 
  assign Queue_17_reset = reset; 
  assign Queue_17_io_enq_valid = _T_180 & _T_144; 
  assign Queue_17_io_enq_bits = auto_in_awuser; 
  assign Queue_17_io_deq_ready = _T_178 & _T_163; 
  assign Queue_18_clock = clock; 
  assign Queue_18_reset = reset; 
  assign Queue_18_io_enq_valid = _T_180 & _T_145; 
  assign Queue_18_io_enq_bits = auto_in_awuser; 
  assign Queue_18_io_deq_ready = _T_178 & _T_164; 
  assign Queue_19_clock = clock; 
  assign Queue_19_reset = reset; 
  assign Queue_19_io_enq_valid = _T_180 & _T_146; 
  assign Queue_19_io_enq_bits = auto_in_awuser; 
  assign Queue_19_io_deq_ready = _T_178 & _T_165; 
  assign Queue_20_clock = clock; 
  assign Queue_20_reset = reset; 
  assign Queue_20_io_enq_valid = _T_180 & _T_147; 
  assign Queue_20_io_enq_bits = auto_in_awuser; 
  assign Queue_20_io_deq_ready = _T_178 & _T_166; 
  assign Queue_21_clock = clock; 
  assign Queue_21_reset = reset; 
  assign Queue_21_io_enq_valid = _T_180 & _T_148; 
  assign Queue_21_io_enq_bits = auto_in_awuser; 
  assign Queue_21_io_deq_ready = _T_178 & _T_167; 
  assign Queue_22_clock = clock; 
  assign Queue_22_reset = reset; 
  assign Queue_22_io_enq_valid = _T_180 & _T_149; 
  assign Queue_22_io_enq_bits = auto_in_awuser; 
  assign Queue_22_io_deq_ready = _T_178 & _T_168; 
  assign Queue_23_clock = clock; 
  assign Queue_23_reset = reset; 
  assign Queue_23_io_enq_valid = _T_180 & _T_150; 
  assign Queue_23_io_enq_bits = auto_in_awuser; 
  assign Queue_23_io_deq_ready = _T_178 & _T_169; 
  assign Queue_24_clock = clock; 
  assign Queue_24_reset = reset; 
  assign Queue_24_io_enq_valid = _T_180 & _T_151; 
  assign Queue_24_io_enq_bits = auto_in_awuser; 
  assign Queue_24_io_deq_ready = _T_178 & _T_170; 
  assign Queue_25_clock = clock; 
  assign Queue_25_reset = reset; 
  assign Queue_25_io_enq_valid = _T_180 & _T_152; 
  assign Queue_25_io_enq_bits = auto_in_awuser; 
  assign Queue_25_io_deq_ready = _T_178 & _T_171; 
  assign Queue_26_clock = clock; 
  assign Queue_26_reset = reset; 
  assign Queue_26_io_enq_valid = _T_180 & _T_153; 
  assign Queue_26_io_enq_bits = auto_in_awuser; 
  assign Queue_26_io_deq_ready = _T_178 & _T_172; 
  assign Queue_27_clock = clock; 
  assign Queue_27_reset = reset; 
  assign Queue_27_io_enq_valid = _T_180 & _T_154; 
  assign Queue_27_io_enq_bits = auto_in_awuser; 
  assign Queue_27_io_deq_ready = _T_178 & _T_173; 
  assign Queue_28_clock = clock; 
  assign Queue_28_reset = reset; 
  assign Queue_28_io_enq_valid = _T_180 & _T_155; 
  assign Queue_28_io_enq_bits = auto_in_awuser; 
  assign Queue_28_io_deq_ready = _T_178 & _T_174; 
  assign Queue_29_clock = clock; 
  assign Queue_29_reset = reset; 
  assign Queue_29_io_enq_valid = _T_180 & _T_156; 
  assign Queue_29_io_enq_bits = auto_in_awuser; 
  assign Queue_29_io_deq_ready = _T_178 & _T_175; 
  assign Queue_30_clock = clock; 
  assign Queue_30_reset = reset; 
  assign Queue_30_io_enq_valid = _T_180 & _T_157; 
  assign Queue_30_io_enq_bits = auto_in_awuser; 
  assign Queue_30_io_deq_ready = _T_178 & _T_176; 
  assign Queue_31_clock = clock; 
  assign Queue_31_reset = reset; 
  assign Queue_31_io_enq_valid = _T_180 & _T_158; 
  assign Queue_31_io_enq_bits = auto_in_awuser; 
  assign Queue_31_io_deq_ready = _T_178 & _T_177; 
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_11) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:54 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_11) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_139) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:75 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_139) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_CAM_9( 
  input         clock, 
  input         reset, 
  output        io_alloc_ready, 
  input         io_alloc_valid, 
  input  [15:0] io_alloc_bits, 
  output [4:0]  io_key, 
  output [15:0] io_data 
);
  reg [15:0] data [0:31]; 
  reg [31:0] _RAND_0;
  wire [15:0] data__T_44_data; 
  wire [4:0] data__T_44_addr; 
  wire [15:0] data__T_41_data; 
  wire [4:0] data__T_41_addr; 
  wire  data__T_41_mask; 
  wire  data__T_41_en; 
  reg [31:0] free; 
  reg [31:0] _RAND_1;
  wire [32:0] _T; 
  wire [31:0] _T_1; 
  wire [31:0] _T_2; 
  wire [33:0] _T_3; 
  wire [31:0] _T_4; 
  wire [31:0] _T_5; 
  wire [35:0] _T_6; 
  wire [31:0] _T_7; 
  wire [31:0] _T_8; 
  wire [39:0] _T_9; 
  wire [31:0] _T_10; 
  wire [31:0] _T_11; 
  wire [47:0] _T_12; 
  wire [31:0] _T_13; 
  wire [31:0] _T_14; 
  wire [32:0] _T_16; 
  wire [32:0] _T_17; 
  wire [32:0] _GEN_11; 
  wire [32:0] free_sel; 
  wire [15:0] _T_18; 
  wire [15:0] _T_19; 
  wire  _T_20; 
  wire [15:0] _T_21; 
  wire [7:0] _T_22; 
  wire [7:0] _T_23; 
  wire  _T_24; 
  wire [7:0] _T_25; 
  wire [3:0] _T_26; 
  wire [3:0] _T_27; 
  wire  _T_28; 
  wire [3:0] _T_29; 
  wire [1:0] _T_30; 
  wire [1:0] _T_31; 
  wire  _T_32; 
  wire [1:0] _T_33; 
  wire  _T_34; 
  wire [3:0] _T_37; 
  wire  _T_40; 
  wire  _T_43; 
  wire  bypass; 
  wire [32:0] clr; 
  wire [32:0] _T_48; 
  wire [32:0] _T_49; 
  assign data__T_44_addr = 5'h0;
  assign data__T_44_data = data[data__T_44_addr]; 
  assign data__T_41_data = io_alloc_bits;
  assign data__T_41_addr = io_key;
  assign data__T_41_mask = 1'h1;
  assign data__T_41_en = io_alloc_ready & io_alloc_valid;
  assign _T = {free, 1'h0}; 
  assign _T_1 = _T[31:0]; 
  assign _T_2 = free | _T_1; 
  assign _T_3 = {_T_2, 2'h0}; 
  assign _T_4 = _T_3[31:0]; 
  assign _T_5 = _T_2 | _T_4; 
  assign _T_6 = {_T_5, 4'h0}; 
  assign _T_7 = _T_6[31:0]; 
  assign _T_8 = _T_5 | _T_7; 
  assign _T_9 = {_T_8, 8'h0}; 
  assign _T_10 = _T_9[31:0]; 
  assign _T_11 = _T_8 | _T_10; 
  assign _T_12 = {_T_11, 16'h0}; 
  assign _T_13 = _T_12[31:0]; 
  assign _T_14 = _T_11 | _T_13; 
  assign _T_16 = {_T_14, 1'h0}; 
  assign _T_17 = ~ _T_16; 
  assign _GEN_11 = {{1'd0}, free}; 
  assign free_sel = _T_17 & _GEN_11; 
  assign _T_18 = free_sel[31:16]; 
  assign _T_19 = free_sel[15:0]; 
  assign _T_20 = _T_18 != 16'h0; 
  assign _T_21 = _T_18 | _T_19; 
  assign _T_22 = _T_21[15:8]; 
  assign _T_23 = _T_21[7:0]; 
  assign _T_24 = _T_22 != 8'h0; 
  assign _T_25 = _T_22 | _T_23; 
  assign _T_26 = _T_25[7:4]; 
  assign _T_27 = _T_25[3:0]; 
  assign _T_28 = _T_26 != 4'h0; 
  assign _T_29 = _T_26 | _T_27; 
  assign _T_30 = _T_29[3:2]; 
  assign _T_31 = _T_29[1:0]; 
  assign _T_32 = _T_30 != 2'h0; 
  assign _T_33 = _T_30 | _T_31; 
  assign _T_34 = _T_33[1]; 
  assign _T_37 = {_T_24,_T_28,_T_32,_T_34}; 
  assign _T_40 = io_alloc_ready & io_alloc_valid; 
  assign _T_43 = 5'h0 == io_key; 
  assign bypass = _T_40 & _T_43; 
  assign clr = _T_40 ? free_sel : 33'h0; 
  assign _T_48 = ~ clr; 
  assign _T_49 = _GEN_11 & _T_48; 
  assign io_alloc_ready = free != 32'h0; 
  assign io_key = {_T_20,_T_37}; 
  assign io_data = bypass ? io_alloc_bits : data__T_44_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    data[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  free = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(data__T_41_en & data__T_41_mask) begin
      data[data__T_41_addr] <= data__T_41_data; 
    end
    if (reset) begin
      free <= 32'hffffffff;
    end else begin
      free <= _T_49[31:0];
    end
  end
endmodule
module dual_CAM( 
  input         clock, 
  input         reset, 
  output        io_alloc_ready, 
  input         io_alloc_valid, 
  input  [15:0] io_alloc_bits, 
  output [2:0]  io_key, 
  input         io_free_valid, 
  input  [2:0]  io_free_bits, 
  output [15:0] io_data 
);
  reg [15:0] data [0:7]; 
  reg [31:0] _RAND_0;
  wire [15:0] data__T_28_data; 
  wire [2:0] data__T_28_addr; 
  wire [15:0] data__T_25_data; 
  wire [2:0] data__T_25_addr; 
  wire  data__T_25_mask; 
  wire  data__T_25_en; 
  reg [7:0] free; 
  reg [31:0] _RAND_1;
  wire [8:0] _T; 
  wire [7:0] _T_1; 
  wire [7:0] _T_2; 
  wire [9:0] _T_3; 
  wire [7:0] _T_4; 
  wire [7:0] _T_5; 
  wire [11:0] _T_6; 
  wire [7:0] _T_7; 
  wire [7:0] _T_8; 
  wire [8:0] _T_10; 
  wire [8:0] _T_11; 
  wire [8:0] _GEN_11; 
  wire [8:0] free_sel; 
  wire [3:0] _T_12; 
  wire [3:0] _T_13; 
  wire  _T_14; 
  wire [3:0] _T_15; 
  wire [1:0] _T_16; 
  wire [1:0] _T_17; 
  wire  _T_18; 
  wire [1:0] _T_19; 
  wire  _T_20; 
  wire [1:0] _T_21; 
  wire  _T_24; 
  wire  _T_27; 
  wire  bypass; 
  wire [8:0] clr; 
  wire [7:0] _T_31; 
  wire [7:0] set; 
  wire [8:0] _T_32; 
  wire [8:0] _T_33; 
  wire [8:0] _GEN_13; 
  wire [8:0] _T_34; 
  assign data__T_28_addr = io_free_bits;
  assign data__T_28_data = data[data__T_28_addr]; 
  assign data__T_25_data = io_alloc_bits;
  assign data__T_25_addr = io_key;
  assign data__T_25_mask = 1'h1;
  assign data__T_25_en = io_alloc_ready & io_alloc_valid;
  assign _T = {free, 1'h0}; 
  assign _T_1 = _T[7:0]; 
  assign _T_2 = free | _T_1; 
  assign _T_3 = {_T_2, 2'h0}; 
  assign _T_4 = _T_3[7:0]; 
  assign _T_5 = _T_2 | _T_4; 
  assign _T_6 = {_T_5, 4'h0}; 
  assign _T_7 = _T_6[7:0]; 
  assign _T_8 = _T_5 | _T_7; 
  assign _T_10 = {_T_8, 1'h0}; 
  assign _T_11 = ~ _T_10; 
  assign _GEN_11 = {{1'd0}, free}; 
  assign free_sel = _T_11 & _GEN_11; 
  assign _T_12 = free_sel[7:4]; 
  assign _T_13 = free_sel[3:0]; 
  assign _T_14 = _T_12 != 4'h0; 
  assign _T_15 = _T_12 | _T_13; 
  assign _T_16 = _T_15[3:2]; 
  assign _T_17 = _T_15[1:0]; 
  assign _T_18 = _T_16 != 2'h0; 
  assign _T_19 = _T_16 | _T_17; 
  assign _T_20 = _T_19[1]; 
  assign _T_21 = {_T_18,_T_20}; 
  assign _T_24 = io_alloc_ready & io_alloc_valid; 
  assign _T_27 = io_free_bits == io_key; 
  assign bypass = _T_24 & _T_27; 
  assign clr = _T_24 ? free_sel : 9'h0; 
  assign _T_31 = 8'h1 << io_free_bits; 
  assign set = io_free_valid ? _T_31 : 8'h0; 
  assign _T_32 = ~ clr; 
  assign _T_33 = _GEN_11 & _T_32; 
  assign _GEN_13 = {{1'd0}, set}; 
  assign _T_34 = _T_33 | _GEN_13; 
  assign io_alloc_ready = free != 8'h0; 
  assign io_key = {_T_14,_T_21}; 
  assign io_data = bypass ? io_alloc_bits : data__T_28_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    data[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  free = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(data__T_25_en & data__T_25_mask) begin
      data[data__T_25_addr] <= data__T_25_data; 
    end
    if (reset) begin
      free <= 8'hff;
    end else begin
      free <= _T_34[7:0];
    end
  end
endmodule
module ChiplinkTop( 
  input         clock, 
  input         reset, 
  output        fpga_io_c2b_clk, 
  output        fpga_io_c2b_rst, 
  output        fpga_io_c2b_send, 
  output [31:0] fpga_io_c2b_data, 
  input         fpga_io_b2c_clk, 
  input         fpga_io_b2c_rst, 
  input         fpga_io_b2c_send, 
  input  [31:0] fpga_io_b2c_data, 
  input         mem_axi4_0_awready, 
  output        mem_axi4_0_awvalid, 
  output [3:0]  mem_axi4_0_awid, 
  output [31:0] mem_axi4_0_awaddr, 
  output [7:0]  mem_axi4_0_awlen, 
  output [2:0]  mem_axi4_0_awsize, 
  output [1:0]  mem_axi4_0_awburst, 
  output        mem_axi4_0_awlock, 
  output [3:0]  mem_axi4_0_awcache, 
  output [2:0]  mem_axi4_0_awprot, 
  output [3:0]  mem_axi4_0_awqos, 
  output [63:0] mem_axi4_0_awinstret, 
  input         mem_axi4_0_wready, 
  output        mem_axi4_0_wvalid, 
  output [63:0] mem_axi4_0_wdata, 
  output [7:0]  mem_axi4_0_wstrb, 
  output        mem_axi4_0_wlast, 
  output        mem_axi4_0_bready, 
  input         mem_axi4_0_bvalid, 
  input  [3:0]  mem_axi4_0_bid, 
  input  [1:0]  mem_axi4_0_bresp, 
  input         mem_axi4_0_arready, 
  output        mem_axi4_0_arvalid, 
  output [3:0]  mem_axi4_0_arid, 
  output [31:0] mem_axi4_0_araddr, 
  output [7:0]  mem_axi4_0_arlen, 
  output [2:0]  mem_axi4_0_arsize, 
  output [1:0]  mem_axi4_0_arburst, 
  output        mem_axi4_0_arlock, 
  output [3:0]  mem_axi4_0_arcache, 
  output [2:0]  mem_axi4_0_arprot, 
  output [3:0]  mem_axi4_0_arqos, 
  output [63:0] mem_axi4_0_arinstret, 
  output        mem_axi4_0_rready, 
  input         mem_axi4_0_rvalid, 
  input  [3:0]  mem_axi4_0_rid, 
  input  [63:0] mem_axi4_0_rdata, 
  input  [1:0]  mem_axi4_0_rresp, 
  input         mem_axi4_0_rlast, 
  input         mmio_axi4_0_awready, 
  output        mmio_axi4_0_awvalid, 
  output        mmio_axi4_0_awid, 
  output [30:0] mmio_axi4_0_awaddr, 
  output [7:0]  mmio_axi4_0_awlen, 
  output [2:0]  mmio_axi4_0_awsize, 
  output [1:0]  mmio_axi4_0_awburst, 
  output        mmio_axi4_0_awlock, 
  output [3:0]  mmio_axi4_0_awcache, 
  output [2:0]  mmio_axi4_0_awprot, 
  output [3:0]  mmio_axi4_0_awqos, 
  output [63:0] mmio_axi4_0_awinstret, 
  input         mmio_axi4_0_wready, 
  output        mmio_axi4_0_wvalid, 
  output [63:0] mmio_axi4_0_wdata, 
  output [7:0]  mmio_axi4_0_wstrb, 
  output        mmio_axi4_0_wlast, 
  output        mmio_axi4_0_bready, 
  input         mmio_axi4_0_bvalid, 
  input  [1:0]  mmio_axi4_0_bresp, 
  input         mmio_axi4_0_arready, 
  output        mmio_axi4_0_arvalid, 
  output        mmio_axi4_0_arid, 
  output [30:0] mmio_axi4_0_araddr, 
  output [7:0]  mmio_axi4_0_arlen, 
  output [2:0]  mmio_axi4_0_arsize, 
  output [1:0]  mmio_axi4_0_arburst, 
  output        mmio_axi4_0_arlock, 
  output [3:0]  mmio_axi4_0_arcache, 
  output [2:0]  mmio_axi4_0_arprot, 
  output [3:0]  mmio_axi4_0_arqos, 
  output [63:0] mmio_axi4_0_arinstret, 
  output        mmio_axi4_0_rready, 
  input         mmio_axi4_0_rvalid, 
  input  [63:0] mmio_axi4_0_rdata, 
  input  [1:0]  mmio_axi4_0_rresp, 
  input         mmio_axi4_0_rlast, 
  output        l2_frontend_bus_axi4_0_awready, 
  input         l2_frontend_bus_axi4_0_awvalid, 
  input  [16:0] l2_frontend_bus_axi4_0_awid, 
  input  [31:0] l2_frontend_bus_axi4_0_awaddr, 
  input  [7:0]  l2_frontend_bus_axi4_0_awlen, 
  input  [2:0]  l2_frontend_bus_axi4_0_awsize, 
  input  [1:0]  l2_frontend_bus_axi4_0_awburst, 
  output        l2_frontend_bus_axi4_0_wready, 
  input         l2_frontend_bus_axi4_0_wvalid, 
  input  [63:0] l2_frontend_bus_axi4_0_wdata, 
  input  [7:0]  l2_frontend_bus_axi4_0_wstrb, 
  input         l2_frontend_bus_axi4_0_wlast, 
  input         l2_frontend_bus_axi4_0_bready, 
  output        l2_frontend_bus_axi4_0_bvalid, 
  output [16:0] l2_frontend_bus_axi4_0_bid, 
  output [1:0]  l2_frontend_bus_axi4_0_bresp, 
  output        l2_frontend_bus_axi4_0_arready, 
  input         l2_frontend_bus_axi4_0_arvalid, 
  input  [16:0] l2_frontend_bus_axi4_0_arid, 
  input  [31:0] l2_frontend_bus_axi4_0_araddr, 
  input  [7:0]  l2_frontend_bus_axi4_0_arlen, 
  input  [2:0]  l2_frontend_bus_axi4_0_arsize, 
  input  [1:0]  l2_frontend_bus_axi4_0_arburst, 
  input         l2_frontend_bus_axi4_0_rready, 
  output        l2_frontend_bus_axi4_0_rvalid, 
  output [16:0] l2_frontend_bus_axi4_0_rid, 
  output [63:0] l2_frontend_bus_axi4_0_rdata, 
  output [1:0]  l2_frontend_bus_axi4_0_rresp, 
  output        l2_frontend_bus_axi4_0_rlast 
);
  wire  xbar_clock; 
  wire  xbar_reset; 
  wire  xbar_auto_in_a_ready; 
  wire  xbar_auto_in_a_valid; 
  wire [2:0] xbar_auto_in_a_bits_opcode; 
  wire [2:0] xbar_auto_in_a_bits_param; 
  wire [3:0] xbar_auto_in_a_bits_size; 
  wire [6:0] xbar_auto_in_a_bits_source; 
  wire [31:0] xbar_auto_in_a_bits_address; 
  wire [7:0] xbar_auto_in_a_bits_mask; 
  wire [63:0] xbar_auto_in_a_bits_data; 
  wire  xbar_auto_in_a_bits_corrupt; 
  wire  xbar_auto_in_c_ready; 
  wire  xbar_auto_in_c_valid; 
  wire [2:0] xbar_auto_in_c_bits_opcode; 
  wire [2:0] xbar_auto_in_c_bits_param; 
  wire [3:0] xbar_auto_in_c_bits_size; 
  wire [6:0] xbar_auto_in_c_bits_source; 
  wire [31:0] xbar_auto_in_c_bits_address; 
  wire  xbar_auto_in_c_bits_corrupt; 
  wire  xbar_auto_in_d_ready; 
  wire  xbar_auto_in_d_valid; 
  wire [2:0] xbar_auto_in_d_bits_opcode; 
  wire [1:0] xbar_auto_in_d_bits_param; 
  wire [3:0] xbar_auto_in_d_bits_size; 
  wire [6:0] xbar_auto_in_d_bits_source; 
  wire  xbar_auto_in_d_bits_sink; 
  wire  xbar_auto_in_d_bits_denied; 
  wire [63:0] xbar_auto_in_d_bits_data; 
  wire  xbar_auto_in_d_bits_corrupt; 
  wire  xbar_auto_in_e_ready; 
  wire  xbar_auto_in_e_valid; 
  wire  xbar_auto_in_e_bits_sink; 
  wire  xbar_auto_out_2_a_ready; 
  wire  xbar_auto_out_2_a_valid; 
  wire [2:0] xbar_auto_out_2_a_bits_opcode; 
  wire [2:0] xbar_auto_out_2_a_bits_param; 
  wire [2:0] xbar_auto_out_2_a_bits_size; 
  wire [6:0] xbar_auto_out_2_a_bits_source; 
  wire [28:0] xbar_auto_out_2_a_bits_address; 
  wire [7:0] xbar_auto_out_2_a_bits_mask; 
  wire  xbar_auto_out_2_a_bits_corrupt; 
  wire  xbar_auto_out_2_c_ready; 
  wire  xbar_auto_out_2_c_valid; 
  wire [2:0] xbar_auto_out_2_c_bits_opcode; 
  wire [2:0] xbar_auto_out_2_c_bits_param; 
  wire [2:0] xbar_auto_out_2_c_bits_size; 
  wire [6:0] xbar_auto_out_2_c_bits_source; 
  wire [28:0] xbar_auto_out_2_c_bits_address; 
  wire  xbar_auto_out_2_c_bits_corrupt; 
  wire  xbar_auto_out_2_d_ready; 
  wire  xbar_auto_out_2_d_valid; 
  wire [2:0] xbar_auto_out_2_d_bits_opcode; 
  wire [1:0] xbar_auto_out_2_d_bits_param; 
  wire [2:0] xbar_auto_out_2_d_bits_size; 
  wire [6:0] xbar_auto_out_2_d_bits_source; 
  wire  xbar_auto_out_2_d_bits_sink; 
  wire  xbar_auto_out_2_d_bits_denied; 
  wire [63:0] xbar_auto_out_2_d_bits_data; 
  wire  xbar_auto_out_2_d_bits_corrupt; 
  wire  xbar_auto_out_2_e_valid; 
  wire  xbar_auto_out_1_a_ready; 
  wire  xbar_auto_out_1_a_valid; 
  wire [2:0] xbar_auto_out_1_a_bits_opcode; 
  wire [2:0] xbar_auto_out_1_a_bits_param; 
  wire [3:0] xbar_auto_out_1_a_bits_size; 
  wire [6:0] xbar_auto_out_1_a_bits_source; 
  wire [30:0] xbar_auto_out_1_a_bits_address; 
  wire [7:0] xbar_auto_out_1_a_bits_mask; 
  wire [63:0] xbar_auto_out_1_a_bits_data; 
  wire  xbar_auto_out_1_a_bits_corrupt; 
  wire  xbar_auto_out_1_d_ready; 
  wire  xbar_auto_out_1_d_valid; 
  wire [2:0] xbar_auto_out_1_d_bits_opcode; 
  wire [3:0] xbar_auto_out_1_d_bits_size; 
  wire [6:0] xbar_auto_out_1_d_bits_source; 
  wire  xbar_auto_out_1_d_bits_denied; 
  wire [63:0] xbar_auto_out_1_d_bits_data; 
  wire  xbar_auto_out_1_d_bits_corrupt; 
  wire  xbar_auto_out_0_a_ready; 
  wire  xbar_auto_out_0_a_valid; 
  wire [2:0] xbar_auto_out_0_a_bits_opcode; 
  wire [2:0] xbar_auto_out_0_a_bits_param; 
  wire [2:0] xbar_auto_out_0_a_bits_size; 
  wire [6:0] xbar_auto_out_0_a_bits_source; 
  wire [31:0] xbar_auto_out_0_a_bits_address; 
  wire [7:0] xbar_auto_out_0_a_bits_mask; 
  wire [63:0] xbar_auto_out_0_a_bits_data; 
  wire  xbar_auto_out_0_a_bits_corrupt; 
  wire  xbar_auto_out_0_d_ready; 
  wire  xbar_auto_out_0_d_valid; 
  wire [2:0] xbar_auto_out_0_d_bits_opcode; 
  wire [2:0] xbar_auto_out_0_d_bits_size; 
  wire [6:0] xbar_auto_out_0_d_bits_source; 
  wire  xbar_auto_out_0_d_bits_denied; 
  wire [63:0] xbar_auto_out_0_d_bits_data; 
  wire  xbar_auto_out_0_d_bits_corrupt; 
  wire  xbar_1_clock; 
  wire  xbar_1_reset; 
  wire  xbar_1_auto_in_a_ready; 
  wire  xbar_1_auto_in_a_valid; 
  wire [2:0] xbar_1_auto_in_a_bits_opcode; 
  wire [2:0] xbar_1_auto_in_a_bits_param; 
  wire [2:0] xbar_1_auto_in_a_bits_size; 
  wire [2:0] xbar_1_auto_in_a_bits_source; 
  wire [31:0] xbar_1_auto_in_a_bits_address; 
  wire [3:0] xbar_1_auto_in_a_bits_mask; 
  wire [31:0] xbar_1_auto_in_a_bits_data; 
  wire  xbar_1_auto_in_a_bits_corrupt; 
  wire  xbar_1_auto_in_d_ready; 
  wire  xbar_1_auto_in_d_valid; 
  wire [2:0] xbar_1_auto_in_d_bits_opcode; 
  wire [1:0] xbar_1_auto_in_d_bits_param; 
  wire [2:0] xbar_1_auto_in_d_bits_size; 
  wire [2:0] xbar_1_auto_in_d_bits_source; 
  wire [5:0] xbar_1_auto_in_d_bits_sink; 
  wire  xbar_1_auto_in_d_bits_denied; 
  wire [31:0] xbar_1_auto_in_d_bits_data; 
  wire  xbar_1_auto_in_d_bits_corrupt; 
  wire  xbar_1_auto_out_1_a_ready; 
  wire  xbar_1_auto_out_1_a_valid; 
  wire [2:0] xbar_1_auto_out_1_a_bits_opcode; 
  wire [2:0] xbar_1_auto_out_1_a_bits_param; 
  wire [2:0] xbar_1_auto_out_1_a_bits_size; 
  wire [2:0] xbar_1_auto_out_1_a_bits_source; 
  wire [28:0] xbar_1_auto_out_1_a_bits_address; 
  wire [3:0] xbar_1_auto_out_1_a_bits_mask; 
  wire  xbar_1_auto_out_1_a_bits_corrupt; 
  wire  xbar_1_auto_out_1_d_ready; 
  wire  xbar_1_auto_out_1_d_valid; 
  wire [2:0] xbar_1_auto_out_1_d_bits_opcode; 
  wire [1:0] xbar_1_auto_out_1_d_bits_param; 
  wire [2:0] xbar_1_auto_out_1_d_bits_size; 
  wire [2:0] xbar_1_auto_out_1_d_bits_source; 
  wire  xbar_1_auto_out_1_d_bits_sink; 
  wire  xbar_1_auto_out_1_d_bits_denied; 
  wire [31:0] xbar_1_auto_out_1_d_bits_data; 
  wire  xbar_1_auto_out_1_d_bits_corrupt; 
  wire  xbar_1_auto_out_0_a_ready; 
  wire  xbar_1_auto_out_0_a_valid; 
  wire [2:0] xbar_1_auto_out_0_a_bits_opcode; 
  wire [2:0] xbar_1_auto_out_0_a_bits_param; 
  wire [2:0] xbar_1_auto_out_0_a_bits_size; 
  wire [2:0] xbar_1_auto_out_0_a_bits_source; 
  wire [31:0] xbar_1_auto_out_0_a_bits_address; 
  wire [3:0] xbar_1_auto_out_0_a_bits_mask; 
  wire [31:0] xbar_1_auto_out_0_a_bits_data; 
  wire  xbar_1_auto_out_0_a_bits_corrupt; 
  wire  xbar_1_auto_out_0_d_ready; 
  wire  xbar_1_auto_out_0_d_valid; 
  wire [2:0] xbar_1_auto_out_0_d_bits_opcode; 
  wire [1:0] xbar_1_auto_out_0_d_bits_param; 
  wire [2:0] xbar_1_auto_out_0_d_bits_size; 
  wire [2:0] xbar_1_auto_out_0_d_bits_source; 
  wire [4:0] xbar_1_auto_out_0_d_bits_sink; 
  wire  xbar_1_auto_out_0_d_bits_denied; 
  wire [31:0] xbar_1_auto_out_0_d_bits_data; 
  wire  xbar_1_auto_out_0_d_bits_corrupt; 
  wire  ferr_clock; 
  wire  ferr_reset; 
  wire  ferr_auto_in_a_ready; 
  wire  ferr_auto_in_a_valid; 
  wire [2:0] ferr_auto_in_a_bits_opcode; 
  wire [2:0] ferr_auto_in_a_bits_param; 
  wire [2:0] ferr_auto_in_a_bits_size; 
  wire [2:0] ferr_auto_in_a_bits_source; 
  wire [28:0] ferr_auto_in_a_bits_address; 
  wire [3:0] ferr_auto_in_a_bits_mask; 
  wire  ferr_auto_in_a_bits_corrupt; 
  wire  ferr_auto_in_d_ready; 
  wire  ferr_auto_in_d_valid; 
  wire [2:0] ferr_auto_in_d_bits_opcode; 
  wire [1:0] ferr_auto_in_d_bits_param; 
  wire [2:0] ferr_auto_in_d_bits_size; 
  wire [2:0] ferr_auto_in_d_bits_source; 
  wire  ferr_auto_in_d_bits_sink; 
  wire  ferr_auto_in_d_bits_denied; 
  wire [31:0] ferr_auto_in_d_bits_data; 
  wire  ferr_auto_in_d_bits_corrupt; 
  wire  chiplink_clock; 
  wire  chiplink_reset; 
  wire  chiplink_auto_mbypass_out_a_ready; 
  wire  chiplink_auto_mbypass_out_a_valid; 
  wire [2:0] chiplink_auto_mbypass_out_a_bits_opcode; 
  wire [2:0] chiplink_auto_mbypass_out_a_bits_param; 
  wire [3:0] chiplink_auto_mbypass_out_a_bits_size; 
  wire [5:0] chiplink_auto_mbypass_out_a_bits_source; 
  wire [31:0] chiplink_auto_mbypass_out_a_bits_address; 
  wire [3:0] chiplink_auto_mbypass_out_a_bits_mask; 
  wire [31:0] chiplink_auto_mbypass_out_a_bits_data; 
  wire  chiplink_auto_mbypass_out_c_ready; 
  wire  chiplink_auto_mbypass_out_c_valid; 
  wire [2:0] chiplink_auto_mbypass_out_c_bits_opcode; 
  wire [2:0] chiplink_auto_mbypass_out_c_bits_param; 
  wire [3:0] chiplink_auto_mbypass_out_c_bits_size; 
  wire [5:0] chiplink_auto_mbypass_out_c_bits_source; 
  wire [31:0] chiplink_auto_mbypass_out_c_bits_address; 
  wire  chiplink_auto_mbypass_out_c_bits_corrupt; 
  wire  chiplink_auto_mbypass_out_d_ready; 
  wire  chiplink_auto_mbypass_out_d_valid; 
  wire [2:0] chiplink_auto_mbypass_out_d_bits_opcode; 
  wire [1:0] chiplink_auto_mbypass_out_d_bits_param; 
  wire [3:0] chiplink_auto_mbypass_out_d_bits_size; 
  wire [5:0] chiplink_auto_mbypass_out_d_bits_source; 
  wire  chiplink_auto_mbypass_out_d_bits_sink; 
  wire  chiplink_auto_mbypass_out_d_bits_denied; 
  wire [31:0] chiplink_auto_mbypass_out_d_bits_data; 
  wire  chiplink_auto_mbypass_out_d_bits_corrupt; 
  wire  chiplink_auto_mbypass_out_e_ready; 
  wire  chiplink_auto_mbypass_out_e_valid; 
  wire  chiplink_auto_mbypass_out_e_bits_sink; 
  wire  chiplink_auto_sbypass_node_in_in_a_ready; 
  wire  chiplink_auto_sbypass_node_in_in_a_valid; 
  wire [2:0] chiplink_auto_sbypass_node_in_in_a_bits_opcode; 
  wire [2:0] chiplink_auto_sbypass_node_in_in_a_bits_param; 
  wire [2:0] chiplink_auto_sbypass_node_in_in_a_bits_size; 
  wire [2:0] chiplink_auto_sbypass_node_in_in_a_bits_source; 
  wire [31:0] chiplink_auto_sbypass_node_in_in_a_bits_address; 
  wire [3:0] chiplink_auto_sbypass_node_in_in_a_bits_mask; 
  wire [31:0] chiplink_auto_sbypass_node_in_in_a_bits_data; 
  wire  chiplink_auto_sbypass_node_in_in_a_bits_corrupt; 
  wire  chiplink_auto_sbypass_node_in_in_d_ready; 
  wire  chiplink_auto_sbypass_node_in_in_d_valid; 
  wire [2:0] chiplink_auto_sbypass_node_in_in_d_bits_opcode; 
  wire [1:0] chiplink_auto_sbypass_node_in_in_d_bits_param; 
  wire [2:0] chiplink_auto_sbypass_node_in_in_d_bits_size; 
  wire [2:0] chiplink_auto_sbypass_node_in_in_d_bits_source; 
  wire [4:0] chiplink_auto_sbypass_node_in_in_d_bits_sink; 
  wire  chiplink_auto_sbypass_node_in_in_d_bits_denied; 
  wire [31:0] chiplink_auto_sbypass_node_in_in_d_bits_data; 
  wire  chiplink_auto_sbypass_node_in_in_d_bits_corrupt; 
  wire  chiplink_auto_io_out_c2b_clk; 
  wire  chiplink_auto_io_out_c2b_rst; 
  wire  chiplink_auto_io_out_c2b_send; 
  wire [31:0] chiplink_auto_io_out_c2b_data; 
  wire  chiplink_auto_io_out_b2c_clk; 
  wire  chiplink_auto_io_out_b2c_rst; 
  wire  chiplink_auto_io_out_b2c_send; 
  wire [31:0] chiplink_auto_io_out_b2c_data; 
  wire  axi4yank_clock; 
  wire  axi4yank_reset; 
  wire  axi4yank_auto_in_awready; 
  wire  axi4yank_auto_in_awvalid; 
  wire [3:0] axi4yank_auto_in_awid; 
  wire [31:0] axi4yank_auto_in_awaddr; 
  wire [7:0] axi4yank_auto_in_awlen; 
  wire [2:0] axi4yank_auto_in_awsize; 
  wire [1:0] axi4yank_auto_in_awburst; 
  wire  axi4yank_auto_in_awlock; 
  wire [3:0] axi4yank_auto_in_awcache; 
  wire [2:0] axi4yank_auto_in_awprot; 
  wire [3:0] axi4yank_auto_in_awqos; 
  wire [11:0] axi4yank_auto_in_awuser; 
  wire [63:0] axi4yank_auto_in_awinstret; 
  wire  axi4yank_auto_in_wready; 
  wire  axi4yank_auto_in_wvalid; 
  wire [63:0] axi4yank_auto_in_wdata; 
  wire [7:0] axi4yank_auto_in_wstrb; 
  wire  axi4yank_auto_in_wlast; 
  wire  axi4yank_auto_in_bready; 
  wire  axi4yank_auto_in_bvalid; 
  wire [3:0] axi4yank_auto_in_bid; 
  wire [1:0] axi4yank_auto_in_bresp; 
  wire [11:0] axi4yank_auto_in_buser; 
  wire  axi4yank_auto_in_arready; 
  wire  axi4yank_auto_in_arvalid; 
  wire [3:0] axi4yank_auto_in_arid; 
  wire [31:0] axi4yank_auto_in_araddr; 
  wire [7:0] axi4yank_auto_in_arlen; 
  wire [2:0] axi4yank_auto_in_arsize; 
  wire [1:0] axi4yank_auto_in_arburst; 
  wire  axi4yank_auto_in_arlock; 
  wire [3:0] axi4yank_auto_in_arcache; 
  wire [2:0] axi4yank_auto_in_arprot; 
  wire [3:0] axi4yank_auto_in_arqos; 
  wire [11:0] axi4yank_auto_in_aruser; 
  wire [63:0] axi4yank_auto_in_arinstret; 
  wire  axi4yank_auto_in_rready; 
  wire  axi4yank_auto_in_rvalid; 
  wire [3:0] axi4yank_auto_in_rid; 
  wire [63:0] axi4yank_auto_in_rdata; 
  wire [1:0] axi4yank_auto_in_rresp; 
  wire [11:0] axi4yank_auto_in_ruser; 
  wire  axi4yank_auto_in_rlast; 
  wire  axi4yank_auto_out_awready; 
  wire  axi4yank_auto_out_awvalid; 
  wire [3:0] axi4yank_auto_out_awid; 
  wire [31:0] axi4yank_auto_out_awaddr; 
  wire [7:0] axi4yank_auto_out_awlen; 
  wire [2:0] axi4yank_auto_out_awsize; 
  wire [1:0] axi4yank_auto_out_awburst; 
  wire  axi4yank_auto_out_awlock; 
  wire [3:0] axi4yank_auto_out_awcache; 
  wire [2:0] axi4yank_auto_out_awprot; 
  wire [3:0] axi4yank_auto_out_awqos; 
  wire [63:0] axi4yank_auto_out_awinstret; 
  wire  axi4yank_auto_out_wready; 
  wire  axi4yank_auto_out_wvalid; 
  wire [63:0] axi4yank_auto_out_wdata; 
  wire [7:0] axi4yank_auto_out_wstrb; 
  wire  axi4yank_auto_out_wlast; 
  wire  axi4yank_auto_out_bready; 
  wire  axi4yank_auto_out_bvalid; 
  wire [3:0] axi4yank_auto_out_bid; 
  wire [1:0] axi4yank_auto_out_bresp; 
  wire  axi4yank_auto_out_arready; 
  wire  axi4yank_auto_out_arvalid; 
  wire [3:0] axi4yank_auto_out_arid; 
  wire [31:0] axi4yank_auto_out_araddr; 
  wire [7:0] axi4yank_auto_out_arlen; 
  wire [2:0] axi4yank_auto_out_arsize; 
  wire [1:0] axi4yank_auto_out_arburst; 
  wire  axi4yank_auto_out_arlock; 
  wire [3:0] axi4yank_auto_out_arcache; 
  wire [2:0] axi4yank_auto_out_arprot; 
  wire [3:0] axi4yank_auto_out_arqos; 
  wire [63:0] axi4yank_auto_out_arinstret; 
  wire  axi4yank_auto_out_rready; 
  wire  axi4yank_auto_out_rvalid; 
  wire [3:0] axi4yank_auto_out_rid; 
  wire [63:0] axi4yank_auto_out_rdata; 
  wire [1:0] axi4yank_auto_out_rresp; 
  wire  axi4yank_auto_out_rlast; 
  wire  axi4index_auto_in_awready; 
  wire  axi4index_auto_in_awvalid; 
  wire [4:0] axi4index_auto_in_awid; 
  wire [31:0] axi4index_auto_in_awaddr; 
  wire [7:0] axi4index_auto_in_awlen; 
  wire [2:0] axi4index_auto_in_awsize; 
  wire [1:0] axi4index_auto_in_awburst; 
  wire  axi4index_auto_in_awlock; 
  wire [3:0] axi4index_auto_in_awcache; 
  wire [2:0] axi4index_auto_in_awprot; 
  wire [3:0] axi4index_auto_in_awqos; 
  wire [10:0] axi4index_auto_in_awuser; 
  wire [63:0] axi4index_auto_in_awinstret; 
  wire  axi4index_auto_in_wready; 
  wire  axi4index_auto_in_wvalid; 
  wire [63:0] axi4index_auto_in_wdata; 
  wire [7:0] axi4index_auto_in_wstrb; 
  wire  axi4index_auto_in_wlast; 
  wire  axi4index_auto_in_bready; 
  wire  axi4index_auto_in_bvalid; 
  wire [4:0] axi4index_auto_in_bid; 
  wire [1:0] axi4index_auto_in_bresp; 
  wire [10:0] axi4index_auto_in_buser; 
  wire  axi4index_auto_in_arready; 
  wire  axi4index_auto_in_arvalid; 
  wire [4:0] axi4index_auto_in_arid; 
  wire [31:0] axi4index_auto_in_araddr; 
  wire [7:0] axi4index_auto_in_arlen; 
  wire [2:0] axi4index_auto_in_arsize; 
  wire [1:0] axi4index_auto_in_arburst; 
  wire  axi4index_auto_in_arlock; 
  wire [3:0] axi4index_auto_in_arcache; 
  wire [2:0] axi4index_auto_in_arprot; 
  wire [3:0] axi4index_auto_in_arqos; 
  wire [10:0] axi4index_auto_in_aruser; 
  wire [63:0] axi4index_auto_in_arinstret; 
  wire  axi4index_auto_in_rready; 
  wire  axi4index_auto_in_rvalid; 
  wire [4:0] axi4index_auto_in_rid; 
  wire [63:0] axi4index_auto_in_rdata; 
  wire [1:0] axi4index_auto_in_rresp; 
  wire [10:0] axi4index_auto_in_ruser; 
  wire  axi4index_auto_in_rlast; 
  wire  axi4index_auto_out_awready; 
  wire  axi4index_auto_out_awvalid; 
  wire [3:0] axi4index_auto_out_awid; 
  wire [31:0] axi4index_auto_out_awaddr; 
  wire [7:0] axi4index_auto_out_awlen; 
  wire [2:0] axi4index_auto_out_awsize; 
  wire [1:0] axi4index_auto_out_awburst; 
  wire  axi4index_auto_out_awlock; 
  wire [3:0] axi4index_auto_out_awcache; 
  wire [2:0] axi4index_auto_out_awprot; 
  wire [3:0] axi4index_auto_out_awqos; 
  wire [11:0] axi4index_auto_out_awuser; 
  wire [63:0] axi4index_auto_out_awinstret; 
  wire  axi4index_auto_out_wready; 
  wire  axi4index_auto_out_wvalid; 
  wire [63:0] axi4index_auto_out_wdata; 
  wire [7:0] axi4index_auto_out_wstrb; 
  wire  axi4index_auto_out_wlast; 
  wire  axi4index_auto_out_bready; 
  wire  axi4index_auto_out_bvalid; 
  wire [3:0] axi4index_auto_out_bid; 
  wire [1:0] axi4index_auto_out_bresp; 
  wire [11:0] axi4index_auto_out_buser; 
  wire  axi4index_auto_out_arready; 
  wire  axi4index_auto_out_arvalid; 
  wire [3:0] axi4index_auto_out_arid; 
  wire [31:0] axi4index_auto_out_araddr; 
  wire [7:0] axi4index_auto_out_arlen; 
  wire [2:0] axi4index_auto_out_arsize; 
  wire [1:0] axi4index_auto_out_arburst; 
  wire  axi4index_auto_out_arlock; 
  wire [3:0] axi4index_auto_out_arcache; 
  wire [2:0] axi4index_auto_out_arprot; 
  wire [3:0] axi4index_auto_out_arqos; 
  wire [11:0] axi4index_auto_out_aruser; 
  wire [63:0] axi4index_auto_out_arinstret; 
  wire  axi4index_auto_out_rready; 
  wire  axi4index_auto_out_rvalid; 
  wire [3:0] axi4index_auto_out_rid; 
  wire [63:0] axi4index_auto_out_rdata; 
  wire [1:0] axi4index_auto_out_rresp; 
  wire [11:0] axi4index_auto_out_ruser; 
  wire  axi4index_auto_out_rlast; 
  wire  tl2axi4_clock; 
  wire  tl2axi4_reset; 
  wire  tl2axi4_auto_in_a_ready; 
  wire  tl2axi4_auto_in_a_valid; 
  wire [2:0] tl2axi4_auto_in_a_bits_opcode; 
  wire [2:0] tl2axi4_auto_in_a_bits_param; 
  wire [2:0] tl2axi4_auto_in_a_bits_size; 
  wire [6:0] tl2axi4_auto_in_a_bits_source; 
  wire [31:0] tl2axi4_auto_in_a_bits_address; 
  wire [7:0] tl2axi4_auto_in_a_bits_mask; 
  wire [63:0] tl2axi4_auto_in_a_bits_data; 
  wire  tl2axi4_auto_in_a_bits_corrupt; 
  wire  tl2axi4_auto_in_d_ready; 
  wire  tl2axi4_auto_in_d_valid; 
  wire [2:0] tl2axi4_auto_in_d_bits_opcode; 
  wire [2:0] tl2axi4_auto_in_d_bits_size; 
  wire [6:0] tl2axi4_auto_in_d_bits_source; 
  wire  tl2axi4_auto_in_d_bits_denied; 
  wire [63:0] tl2axi4_auto_in_d_bits_data; 
  wire  tl2axi4_auto_in_d_bits_corrupt; 
  wire  tl2axi4_auto_out_awready; 
  wire  tl2axi4_auto_out_awvalid; 
  wire [4:0] tl2axi4_auto_out_awid; 
  wire [31:0] tl2axi4_auto_out_awaddr; 
  wire [7:0] tl2axi4_auto_out_awlen; 
  wire [2:0] tl2axi4_auto_out_awsize; 
  wire [1:0] tl2axi4_auto_out_awburst; 
  wire  tl2axi4_auto_out_awlock; 
  wire [3:0] tl2axi4_auto_out_awcache; 
  wire [2:0] tl2axi4_auto_out_awprot; 
  wire [3:0] tl2axi4_auto_out_awqos; 
  wire [10:0] tl2axi4_auto_out_awuser; 
  wire [63:0] tl2axi4_auto_out_awinstret; 
  wire  tl2axi4_auto_out_wready; 
  wire  tl2axi4_auto_out_wvalid; 
  wire [63:0] tl2axi4_auto_out_wdata; 
  wire [7:0] tl2axi4_auto_out_wstrb; 
  wire  tl2axi4_auto_out_wlast; 
  wire  tl2axi4_auto_out_bready; 
  wire  tl2axi4_auto_out_bvalid; 
  wire [4:0] tl2axi4_auto_out_bid; 
  wire [1:0] tl2axi4_auto_out_bresp; 
  wire [10:0] tl2axi4_auto_out_buser; 
  wire  tl2axi4_auto_out_arready; 
  wire  tl2axi4_auto_out_arvalid; 
  wire [4:0] tl2axi4_auto_out_arid; 
  wire [31:0] tl2axi4_auto_out_araddr; 
  wire [7:0] tl2axi4_auto_out_arlen; 
  wire [2:0] tl2axi4_auto_out_arsize; 
  wire [1:0] tl2axi4_auto_out_arburst; 
  wire  tl2axi4_auto_out_arlock; 
  wire [3:0] tl2axi4_auto_out_arcache; 
  wire [2:0] tl2axi4_auto_out_arprot; 
  wire [3:0] tl2axi4_auto_out_arqos; 
  wire [10:0] tl2axi4_auto_out_aruser; 
  wire [63:0] tl2axi4_auto_out_arinstret; 
  wire  tl2axi4_auto_out_rready; 
  wire  tl2axi4_auto_out_rvalid; 
  wire [4:0] tl2axi4_auto_out_rid; 
  wire [63:0] tl2axi4_auto_out_rdata; 
  wire [1:0] tl2axi4_auto_out_rresp; 
  wire [10:0] tl2axi4_auto_out_ruser; 
  wire  tl2axi4_auto_out_rlast; 
  wire  axi4buf_clock; 
  wire  axi4buf_reset; 
  wire  axi4buf_auto_in_awready; 
  wire  axi4buf_auto_in_awvalid; 
  wire [30:0] axi4buf_auto_in_awaddr; 
  wire [7:0] axi4buf_auto_in_awlen; 
  wire [2:0] axi4buf_auto_in_awsize; 
  wire [1:0] axi4buf_auto_in_awburst; 
  wire  axi4buf_auto_in_awlock; 
  wire [3:0] axi4buf_auto_in_awcache; 
  wire [2:0] axi4buf_auto_in_awprot; 
  wire [3:0] axi4buf_auto_in_awqos; 
  wire [63:0] axi4buf_auto_in_awinstret; 
  wire  axi4buf_auto_in_wready; 
  wire  axi4buf_auto_in_wvalid; 
  wire [63:0] axi4buf_auto_in_wdata; 
  wire [7:0] axi4buf_auto_in_wstrb; 
  wire  axi4buf_auto_in_wlast; 
  wire  axi4buf_auto_in_bready; 
  wire  axi4buf_auto_in_bvalid; 
  wire [1:0] axi4buf_auto_in_bresp; 
  wire  axi4buf_auto_in_arready; 
  wire  axi4buf_auto_in_arvalid; 
  wire [30:0] axi4buf_auto_in_araddr; 
  wire [7:0] axi4buf_auto_in_arlen; 
  wire [2:0] axi4buf_auto_in_arsize; 
  wire [1:0] axi4buf_auto_in_arburst; 
  wire  axi4buf_auto_in_arlock; 
  wire [3:0] axi4buf_auto_in_arcache; 
  wire [2:0] axi4buf_auto_in_arprot; 
  wire [3:0] axi4buf_auto_in_arqos; 
  wire [63:0] axi4buf_auto_in_arinstret; 
  wire  axi4buf_auto_in_rready; 
  wire  axi4buf_auto_in_rvalid; 
  wire [63:0] axi4buf_auto_in_rdata; 
  wire [1:0] axi4buf_auto_in_rresp; 
  wire  axi4buf_auto_in_rlast; 
  wire  axi4buf_auto_out_awready; 
  wire  axi4buf_auto_out_awvalid; 
  wire  axi4buf_auto_out_awid; 
  wire [30:0] axi4buf_auto_out_awaddr; 
  wire [7:0] axi4buf_auto_out_awlen; 
  wire [2:0] axi4buf_auto_out_awsize; 
  wire [1:0] axi4buf_auto_out_awburst; 
  wire  axi4buf_auto_out_awlock; 
  wire [3:0] axi4buf_auto_out_awcache; 
  wire [2:0] axi4buf_auto_out_awprot; 
  wire [3:0] axi4buf_auto_out_awqos; 
  wire [63:0] axi4buf_auto_out_awinstret; 
  wire  axi4buf_auto_out_wready; 
  wire  axi4buf_auto_out_wvalid; 
  wire [63:0] axi4buf_auto_out_wdata; 
  wire [7:0] axi4buf_auto_out_wstrb; 
  wire  axi4buf_auto_out_wlast; 
  wire  axi4buf_auto_out_bready; 
  wire  axi4buf_auto_out_bvalid; 
  wire [1:0] axi4buf_auto_out_bresp; 
  wire  axi4buf_auto_out_arready; 
  wire  axi4buf_auto_out_arvalid; 
  wire  axi4buf_auto_out_arid; 
  wire [30:0] axi4buf_auto_out_araddr; 
  wire [7:0] axi4buf_auto_out_arlen; 
  wire [2:0] axi4buf_auto_out_arsize; 
  wire [1:0] axi4buf_auto_out_arburst; 
  wire  axi4buf_auto_out_arlock; 
  wire [3:0] axi4buf_auto_out_arcache; 
  wire [2:0] axi4buf_auto_out_arprot; 
  wire [3:0] axi4buf_auto_out_arqos; 
  wire [63:0] axi4buf_auto_out_arinstret; 
  wire  axi4buf_auto_out_rready; 
  wire  axi4buf_auto_out_rvalid; 
  wire [63:0] axi4buf_auto_out_rdata; 
  wire [1:0] axi4buf_auto_out_rresp; 
  wire  axi4buf_auto_out_rlast; 
  wire  axi4yank_1_clock; 
  wire  axi4yank_1_reset; 
  wire  axi4yank_1_auto_in_awready; 
  wire  axi4yank_1_auto_in_awvalid; 
  wire [30:0] axi4yank_1_auto_in_awaddr; 
  wire [7:0] axi4yank_1_auto_in_awlen; 
  wire [2:0] axi4yank_1_auto_in_awsize; 
  wire [1:0] axi4yank_1_auto_in_awburst; 
  wire  axi4yank_1_auto_in_awlock; 
  wire [3:0] axi4yank_1_auto_in_awcache; 
  wire [2:0] axi4yank_1_auto_in_awprot; 
  wire [3:0] axi4yank_1_auto_in_awqos; 
  wire [15:0] axi4yank_1_auto_in_awuser; 
  wire [63:0] axi4yank_1_auto_in_awinstret; 
  wire  axi4yank_1_auto_in_wready; 
  wire  axi4yank_1_auto_in_wvalid; 
  wire [63:0] axi4yank_1_auto_in_wdata; 
  wire [7:0] axi4yank_1_auto_in_wstrb; 
  wire  axi4yank_1_auto_in_wlast; 
  wire  axi4yank_1_auto_in_bready; 
  wire  axi4yank_1_auto_in_bvalid; 
  wire [1:0] axi4yank_1_auto_in_bresp; 
  wire [15:0] axi4yank_1_auto_in_buser; 
  wire  axi4yank_1_auto_in_arready; 
  wire  axi4yank_1_auto_in_arvalid; 
  wire [30:0] axi4yank_1_auto_in_araddr; 
  wire [7:0] axi4yank_1_auto_in_arlen; 
  wire [2:0] axi4yank_1_auto_in_arsize; 
  wire [1:0] axi4yank_1_auto_in_arburst; 
  wire  axi4yank_1_auto_in_arlock; 
  wire [3:0] axi4yank_1_auto_in_arcache; 
  wire [2:0] axi4yank_1_auto_in_arprot; 
  wire [3:0] axi4yank_1_auto_in_arqos; 
  wire [15:0] axi4yank_1_auto_in_aruser; 
  wire [63:0] axi4yank_1_auto_in_arinstret; 
  wire  axi4yank_1_auto_in_rready; 
  wire  axi4yank_1_auto_in_rvalid; 
  wire [63:0] axi4yank_1_auto_in_rdata; 
  wire [1:0] axi4yank_1_auto_in_rresp; 
  wire [15:0] axi4yank_1_auto_in_ruser; 
  wire  axi4yank_1_auto_in_rlast; 
  wire  axi4yank_1_auto_out_awready; 
  wire  axi4yank_1_auto_out_awvalid; 
  wire [30:0] axi4yank_1_auto_out_awaddr; 
  wire [7:0] axi4yank_1_auto_out_awlen; 
  wire [2:0] axi4yank_1_auto_out_awsize; 
  wire [1:0] axi4yank_1_auto_out_awburst; 
  wire  axi4yank_1_auto_out_awlock; 
  wire [3:0] axi4yank_1_auto_out_awcache; 
  wire [2:0] axi4yank_1_auto_out_awprot; 
  wire [3:0] axi4yank_1_auto_out_awqos; 
  wire [63:0] axi4yank_1_auto_out_awinstret; 
  wire  axi4yank_1_auto_out_wready; 
  wire  axi4yank_1_auto_out_wvalid; 
  wire [63:0] axi4yank_1_auto_out_wdata; 
  wire [7:0] axi4yank_1_auto_out_wstrb; 
  wire  axi4yank_1_auto_out_wlast; 
  wire  axi4yank_1_auto_out_bready; 
  wire  axi4yank_1_auto_out_bvalid; 
  wire [1:0] axi4yank_1_auto_out_bresp; 
  wire  axi4yank_1_auto_out_arready; 
  wire  axi4yank_1_auto_out_arvalid; 
  wire [30:0] axi4yank_1_auto_out_araddr; 
  wire [7:0] axi4yank_1_auto_out_arlen; 
  wire [2:0] axi4yank_1_auto_out_arsize; 
  wire [1:0] axi4yank_1_auto_out_arburst; 
  wire  axi4yank_1_auto_out_arlock; 
  wire [3:0] axi4yank_1_auto_out_arcache; 
  wire [2:0] axi4yank_1_auto_out_arprot; 
  wire [3:0] axi4yank_1_auto_out_arqos; 
  wire [63:0] axi4yank_1_auto_out_arinstret; 
  wire  axi4yank_1_auto_out_rready; 
  wire  axi4yank_1_auto_out_rvalid; 
  wire [63:0] axi4yank_1_auto_out_rdata; 
  wire [1:0] axi4yank_1_auto_out_rresp; 
  wire  axi4yank_1_auto_out_rlast; 
  wire  axi4deint_clock; 
  wire  axi4deint_reset; 
  wire  axi4deint_auto_in_awready; 
  wire  axi4deint_auto_in_awvalid; 
  wire [30:0] axi4deint_auto_in_awaddr; 
  wire [7:0] axi4deint_auto_in_awlen; 
  wire [2:0] axi4deint_auto_in_awsize; 
  wire [1:0] axi4deint_auto_in_awburst; 
  wire  axi4deint_auto_in_awlock; 
  wire [3:0] axi4deint_auto_in_awcache; 
  wire [2:0] axi4deint_auto_in_awprot; 
  wire [3:0] axi4deint_auto_in_awqos; 
  wire [15:0] axi4deint_auto_in_awuser; 
  wire [63:0] axi4deint_auto_in_awinstret; 
  wire  axi4deint_auto_in_wready; 
  wire  axi4deint_auto_in_wvalid; 
  wire [63:0] axi4deint_auto_in_wdata; 
  wire [7:0] axi4deint_auto_in_wstrb; 
  wire  axi4deint_auto_in_wlast; 
  wire  axi4deint_auto_in_bready; 
  wire  axi4deint_auto_in_bvalid; 
  wire [1:0] axi4deint_auto_in_bresp; 
  wire [15:0] axi4deint_auto_in_buser; 
  wire  axi4deint_auto_in_arready; 
  wire  axi4deint_auto_in_arvalid; 
  wire [30:0] axi4deint_auto_in_araddr; 
  wire [7:0] axi4deint_auto_in_arlen; 
  wire [2:0] axi4deint_auto_in_arsize; 
  wire [1:0] axi4deint_auto_in_arburst; 
  wire  axi4deint_auto_in_arlock; 
  wire [3:0] axi4deint_auto_in_arcache; 
  wire [2:0] axi4deint_auto_in_arprot; 
  wire [3:0] axi4deint_auto_in_arqos; 
  wire [15:0] axi4deint_auto_in_aruser; 
  wire [63:0] axi4deint_auto_in_arinstret; 
  wire  axi4deint_auto_in_rready; 
  wire  axi4deint_auto_in_rvalid; 
  wire [63:0] axi4deint_auto_in_rdata; 
  wire [1:0] axi4deint_auto_in_rresp; 
  wire [15:0] axi4deint_auto_in_ruser; 
  wire  axi4deint_auto_in_rlast; 
  wire  axi4deint_auto_out_awready; 
  wire  axi4deint_auto_out_awvalid; 
  wire [30:0] axi4deint_auto_out_awaddr; 
  wire [7:0] axi4deint_auto_out_awlen; 
  wire [2:0] axi4deint_auto_out_awsize; 
  wire [1:0] axi4deint_auto_out_awburst; 
  wire  axi4deint_auto_out_awlock; 
  wire [3:0] axi4deint_auto_out_awcache; 
  wire [2:0] axi4deint_auto_out_awprot; 
  wire [3:0] axi4deint_auto_out_awqos; 
  wire [15:0] axi4deint_auto_out_awuser; 
  wire [63:0] axi4deint_auto_out_awinstret; 
  wire  axi4deint_auto_out_wready; 
  wire  axi4deint_auto_out_wvalid; 
  wire [63:0] axi4deint_auto_out_wdata; 
  wire [7:0] axi4deint_auto_out_wstrb; 
  wire  axi4deint_auto_out_wlast; 
  wire  axi4deint_auto_out_bready; 
  wire  axi4deint_auto_out_bvalid; 
  wire [1:0] axi4deint_auto_out_bresp; 
  wire [15:0] axi4deint_auto_out_buser; 
  wire  axi4deint_auto_out_arready; 
  wire  axi4deint_auto_out_arvalid; 
  wire [30:0] axi4deint_auto_out_araddr; 
  wire [7:0] axi4deint_auto_out_arlen; 
  wire [2:0] axi4deint_auto_out_arsize; 
  wire [1:0] axi4deint_auto_out_arburst; 
  wire  axi4deint_auto_out_arlock; 
  wire [3:0] axi4deint_auto_out_arcache; 
  wire [2:0] axi4deint_auto_out_arprot; 
  wire [3:0] axi4deint_auto_out_arqos; 
  wire [15:0] axi4deint_auto_out_aruser; 
  wire [63:0] axi4deint_auto_out_arinstret; 
  wire  axi4deint_auto_out_rready; 
  wire  axi4deint_auto_out_rvalid; 
  wire [63:0] axi4deint_auto_out_rdata; 
  wire [1:0] axi4deint_auto_out_rresp; 
  wire [15:0] axi4deint_auto_out_ruser; 
  wire  axi4deint_auto_out_rlast; 
  wire  axi4index_1_auto_in_awready; 
  wire  axi4index_1_auto_in_awvalid; 
  wire [4:0] axi4index_1_auto_in_awid; 
  wire [30:0] axi4index_1_auto_in_awaddr; 
  wire [7:0] axi4index_1_auto_in_awlen; 
  wire [2:0] axi4index_1_auto_in_awsize; 
  wire [1:0] axi4index_1_auto_in_awburst; 
  wire  axi4index_1_auto_in_awlock; 
  wire [3:0] axi4index_1_auto_in_awcache; 
  wire [2:0] axi4index_1_auto_in_awprot; 
  wire [3:0] axi4index_1_auto_in_awqos; 
  wire [10:0] axi4index_1_auto_in_awuser; 
  wire [63:0] axi4index_1_auto_in_awinstret; 
  wire  axi4index_1_auto_in_wready; 
  wire  axi4index_1_auto_in_wvalid; 
  wire [63:0] axi4index_1_auto_in_wdata; 
  wire [7:0] axi4index_1_auto_in_wstrb; 
  wire  axi4index_1_auto_in_wlast; 
  wire  axi4index_1_auto_in_bready; 
  wire  axi4index_1_auto_in_bvalid; 
  wire [4:0] axi4index_1_auto_in_bid; 
  wire [1:0] axi4index_1_auto_in_bresp; 
  wire [10:0] axi4index_1_auto_in_buser; 
  wire  axi4index_1_auto_in_arready; 
  wire  axi4index_1_auto_in_arvalid; 
  wire [4:0] axi4index_1_auto_in_arid; 
  wire [30:0] axi4index_1_auto_in_araddr; 
  wire [7:0] axi4index_1_auto_in_arlen; 
  wire [2:0] axi4index_1_auto_in_arsize; 
  wire [1:0] axi4index_1_auto_in_arburst; 
  wire  axi4index_1_auto_in_arlock; 
  wire [3:0] axi4index_1_auto_in_arcache; 
  wire [2:0] axi4index_1_auto_in_arprot; 
  wire [3:0] axi4index_1_auto_in_arqos; 
  wire [10:0] axi4index_1_auto_in_aruser; 
  wire [63:0] axi4index_1_auto_in_arinstret; 
  wire  axi4index_1_auto_in_rready; 
  wire  axi4index_1_auto_in_rvalid; 
  wire [4:0] axi4index_1_auto_in_rid; 
  wire [63:0] axi4index_1_auto_in_rdata; 
  wire [1:0] axi4index_1_auto_in_rresp; 
  wire [10:0] axi4index_1_auto_in_ruser; 
  wire  axi4index_1_auto_in_rlast; 
  wire  axi4index_1_auto_out_awready; 
  wire  axi4index_1_auto_out_awvalid; 
  wire [30:0] axi4index_1_auto_out_awaddr; 
  wire [7:0] axi4index_1_auto_out_awlen; 
  wire [2:0] axi4index_1_auto_out_awsize; 
  wire [1:0] axi4index_1_auto_out_awburst; 
  wire  axi4index_1_auto_out_awlock; 
  wire [3:0] axi4index_1_auto_out_awcache; 
  wire [2:0] axi4index_1_auto_out_awprot; 
  wire [3:0] axi4index_1_auto_out_awqos; 
  wire [15:0] axi4index_1_auto_out_awuser; 
  wire [63:0] axi4index_1_auto_out_awinstret; 
  wire  axi4index_1_auto_out_wready; 
  wire  axi4index_1_auto_out_wvalid; 
  wire [63:0] axi4index_1_auto_out_wdata; 
  wire [7:0] axi4index_1_auto_out_wstrb; 
  wire  axi4index_1_auto_out_wlast; 
  wire  axi4index_1_auto_out_bready; 
  wire  axi4index_1_auto_out_bvalid; 
  wire [1:0] axi4index_1_auto_out_bresp; 
  wire [15:0] axi4index_1_auto_out_buser; 
  wire  axi4index_1_auto_out_arready; 
  wire  axi4index_1_auto_out_arvalid; 
  wire [30:0] axi4index_1_auto_out_araddr; 
  wire [7:0] axi4index_1_auto_out_arlen; 
  wire [2:0] axi4index_1_auto_out_arsize; 
  wire [1:0] axi4index_1_auto_out_arburst; 
  wire  axi4index_1_auto_out_arlock; 
  wire [3:0] axi4index_1_auto_out_arcache; 
  wire [2:0] axi4index_1_auto_out_arprot; 
  wire [3:0] axi4index_1_auto_out_arqos; 
  wire [15:0] axi4index_1_auto_out_aruser; 
  wire [63:0] axi4index_1_auto_out_arinstret; 
  wire  axi4index_1_auto_out_rready; 
  wire  axi4index_1_auto_out_rvalid; 
  wire [63:0] axi4index_1_auto_out_rdata; 
  wire [1:0] axi4index_1_auto_out_rresp; 
  wire [15:0] axi4index_1_auto_out_ruser; 
  wire  axi4index_1_auto_out_rlast; 
  wire  tl2axi4_1_clock; 
  wire  tl2axi4_1_reset; 
  wire  tl2axi4_1_auto_in_a_ready; 
  wire  tl2axi4_1_auto_in_a_valid; 
  wire [2:0] tl2axi4_1_auto_in_a_bits_opcode; 
  wire [2:0] tl2axi4_1_auto_in_a_bits_param; 
  wire [3:0] tl2axi4_1_auto_in_a_bits_size; 
  wire [6:0] tl2axi4_1_auto_in_a_bits_source; 
  wire [30:0] tl2axi4_1_auto_in_a_bits_address; 
  wire [7:0] tl2axi4_1_auto_in_a_bits_mask; 
  wire [63:0] tl2axi4_1_auto_in_a_bits_data; 
  wire  tl2axi4_1_auto_in_a_bits_corrupt; 
  wire  tl2axi4_1_auto_in_d_ready; 
  wire  tl2axi4_1_auto_in_d_valid; 
  wire [2:0] tl2axi4_1_auto_in_d_bits_opcode; 
  wire [3:0] tl2axi4_1_auto_in_d_bits_size; 
  wire [6:0] tl2axi4_1_auto_in_d_bits_source; 
  wire  tl2axi4_1_auto_in_d_bits_denied; 
  wire [63:0] tl2axi4_1_auto_in_d_bits_data; 
  wire  tl2axi4_1_auto_in_d_bits_corrupt; 
  wire  tl2axi4_1_auto_out_awready; 
  wire  tl2axi4_1_auto_out_awvalid; 
  wire [4:0] tl2axi4_1_auto_out_awid; 
  wire [30:0] tl2axi4_1_auto_out_awaddr; 
  wire [7:0] tl2axi4_1_auto_out_awlen; 
  wire [2:0] tl2axi4_1_auto_out_awsize; 
  wire [1:0] tl2axi4_1_auto_out_awburst; 
  wire  tl2axi4_1_auto_out_awlock; 
  wire [3:0] tl2axi4_1_auto_out_awcache; 
  wire [2:0] tl2axi4_1_auto_out_awprot; 
  wire [3:0] tl2axi4_1_auto_out_awqos; 
  wire [10:0] tl2axi4_1_auto_out_awuser; 
  wire [63:0] tl2axi4_1_auto_out_awinstret; 
  wire  tl2axi4_1_auto_out_wready; 
  wire  tl2axi4_1_auto_out_wvalid; 
  wire [63:0] tl2axi4_1_auto_out_wdata; 
  wire [7:0] tl2axi4_1_auto_out_wstrb; 
  wire  tl2axi4_1_auto_out_wlast; 
  wire  tl2axi4_1_auto_out_bready; 
  wire  tl2axi4_1_auto_out_bvalid; 
  wire [4:0] tl2axi4_1_auto_out_bid; 
  wire [1:0] tl2axi4_1_auto_out_bresp; 
  wire [10:0] tl2axi4_1_auto_out_buser; 
  wire  tl2axi4_1_auto_out_arready; 
  wire  tl2axi4_1_auto_out_arvalid; 
  wire [4:0] tl2axi4_1_auto_out_arid; 
  wire [30:0] tl2axi4_1_auto_out_araddr; 
  wire [7:0] tl2axi4_1_auto_out_arlen; 
  wire [2:0] tl2axi4_1_auto_out_arsize; 
  wire [1:0] tl2axi4_1_auto_out_arburst; 
  wire  tl2axi4_1_auto_out_arlock; 
  wire [3:0] tl2axi4_1_auto_out_arcache; 
  wire [2:0] tl2axi4_1_auto_out_arprot; 
  wire [3:0] tl2axi4_1_auto_out_arqos; 
  wire [10:0] tl2axi4_1_auto_out_aruser; 
  wire [63:0] tl2axi4_1_auto_out_arinstret; 
  wire  tl2axi4_1_auto_out_rready; 
  wire  tl2axi4_1_auto_out_rvalid; 
  wire [4:0] tl2axi4_1_auto_out_rid; 
  wire [63:0] tl2axi4_1_auto_out_rdata; 
  wire [1:0] tl2axi4_1_auto_out_rresp; 
  wire [10:0] tl2axi4_1_auto_out_ruser; 
  wire  tl2axi4_1_auto_out_rlast; 
  wire  fixer_clock; 
  wire  fixer_reset; 
  wire  fixer_auto_in_a_ready; 
  wire  fixer_auto_in_a_valid; 
  wire [2:0] fixer_auto_in_a_bits_opcode; 
  wire [2:0] fixer_auto_in_a_bits_param; 
  wire [2:0] fixer_auto_in_a_bits_size; 
  wire [2:0] fixer_auto_in_a_bits_source; 
  wire [31:0] fixer_auto_in_a_bits_address; 
  wire [3:0] fixer_auto_in_a_bits_mask; 
  wire [31:0] fixer_auto_in_a_bits_data; 
  wire  fixer_auto_in_a_bits_corrupt; 
  wire  fixer_auto_in_d_ready; 
  wire  fixer_auto_in_d_valid; 
  wire [2:0] fixer_auto_in_d_bits_opcode; 
  wire [1:0] fixer_auto_in_d_bits_param; 
  wire [2:0] fixer_auto_in_d_bits_size; 
  wire [2:0] fixer_auto_in_d_bits_source; 
  wire [5:0] fixer_auto_in_d_bits_sink; 
  wire  fixer_auto_in_d_bits_denied; 
  wire [31:0] fixer_auto_in_d_bits_data; 
  wire  fixer_auto_in_d_bits_corrupt; 
  wire  fixer_auto_out_a_ready; 
  wire  fixer_auto_out_a_valid; 
  wire [2:0] fixer_auto_out_a_bits_opcode; 
  wire [2:0] fixer_auto_out_a_bits_param; 
  wire [2:0] fixer_auto_out_a_bits_size; 
  wire [2:0] fixer_auto_out_a_bits_source; 
  wire [31:0] fixer_auto_out_a_bits_address; 
  wire [3:0] fixer_auto_out_a_bits_mask; 
  wire [31:0] fixer_auto_out_a_bits_data; 
  wire  fixer_auto_out_a_bits_corrupt; 
  wire  fixer_auto_out_d_ready; 
  wire  fixer_auto_out_d_valid; 
  wire [2:0] fixer_auto_out_d_bits_opcode; 
  wire [1:0] fixer_auto_out_d_bits_param; 
  wire [2:0] fixer_auto_out_d_bits_size; 
  wire [2:0] fixer_auto_out_d_bits_source; 
  wire [5:0] fixer_auto_out_d_bits_sink; 
  wire  fixer_auto_out_d_bits_denied; 
  wire [31:0] fixer_auto_out_d_bits_data; 
  wire  fixer_auto_out_d_bits_corrupt; 
  wire  widget_clock; 
  wire  widget_reset; 
  wire  widget_auto_in_a_ready; 
  wire  widget_auto_in_a_valid; 
  wire [2:0] widget_auto_in_a_bits_opcode; 
  wire [2:0] widget_auto_in_a_bits_param; 
  wire [2:0] widget_auto_in_a_bits_size; 
  wire [2:0] widget_auto_in_a_bits_source; 
  wire [31:0] widget_auto_in_a_bits_address; 
  wire [7:0] widget_auto_in_a_bits_mask; 
  wire [63:0] widget_auto_in_a_bits_data; 
  wire  widget_auto_in_a_bits_corrupt; 
  wire  widget_auto_in_d_ready; 
  wire  widget_auto_in_d_valid; 
  wire [2:0] widget_auto_in_d_bits_opcode; 
  wire [2:0] widget_auto_in_d_bits_size; 
  wire [2:0] widget_auto_in_d_bits_source; 
  wire  widget_auto_in_d_bits_denied; 
  wire [63:0] widget_auto_in_d_bits_data; 
  wire  widget_auto_in_d_bits_corrupt; 
  wire  widget_auto_out_a_ready; 
  wire  widget_auto_out_a_valid; 
  wire [2:0] widget_auto_out_a_bits_opcode; 
  wire [2:0] widget_auto_out_a_bits_param; 
  wire [2:0] widget_auto_out_a_bits_size; 
  wire [2:0] widget_auto_out_a_bits_source; 
  wire [31:0] widget_auto_out_a_bits_address; 
  wire [3:0] widget_auto_out_a_bits_mask; 
  wire [31:0] widget_auto_out_a_bits_data; 
  wire  widget_auto_out_a_bits_corrupt; 
  wire  widget_auto_out_d_ready; 
  wire  widget_auto_out_d_valid; 
  wire [2:0] widget_auto_out_d_bits_opcode; 
  wire [1:0] widget_auto_out_d_bits_param; 
  wire [2:0] widget_auto_out_d_bits_size; 
  wire [2:0] widget_auto_out_d_bits_source; 
  wire [5:0] widget_auto_out_d_bits_sink; 
  wire  widget_auto_out_d_bits_denied; 
  wire [31:0] widget_auto_out_d_bits_data; 
  wire  widget_auto_out_d_bits_corrupt; 
  wire  axi42tl_clock; 
  wire  axi42tl_reset; 
  wire  axi42tl_auto_in_awready; 
  wire  axi42tl_auto_in_awvalid; 
  wire  axi42tl_auto_in_awid; 
  wire [31:0] axi42tl_auto_in_awaddr; 
  wire [7:0] axi42tl_auto_in_awlen; 
  wire [2:0] axi42tl_auto_in_awsize; 
  wire  axi42tl_auto_in_wready; 
  wire  axi42tl_auto_in_wvalid; 
  wire [63:0] axi42tl_auto_in_wdata; 
  wire [7:0] axi42tl_auto_in_wstrb; 
  wire  axi42tl_auto_in_wlast; 
  wire  axi42tl_auto_in_bready; 
  wire  axi42tl_auto_in_bvalid; 
  wire  axi42tl_auto_in_bid; 
  wire [1:0] axi42tl_auto_in_bresp; 
  wire  axi42tl_auto_in_arready; 
  wire  axi42tl_auto_in_arvalid; 
  wire  axi42tl_auto_in_arid; 
  wire [31:0] axi42tl_auto_in_araddr; 
  wire [7:0] axi42tl_auto_in_arlen; 
  wire [2:0] axi42tl_auto_in_arsize; 
  wire  axi42tl_auto_in_rready; 
  wire  axi42tl_auto_in_rvalid; 
  wire  axi42tl_auto_in_rid; 
  wire [63:0] axi42tl_auto_in_rdata; 
  wire [1:0] axi42tl_auto_in_rresp; 
  wire  axi42tl_auto_in_rlast; 
  wire  axi42tl_auto_out_a_ready; 
  wire  axi42tl_auto_out_a_valid; 
  wire [2:0] axi42tl_auto_out_a_bits_opcode; 
  wire [2:0] axi42tl_auto_out_a_bits_param; 
  wire [2:0] axi42tl_auto_out_a_bits_size; 
  wire [2:0] axi42tl_auto_out_a_bits_source; 
  wire [31:0] axi42tl_auto_out_a_bits_address; 
  wire [7:0] axi42tl_auto_out_a_bits_mask; 
  wire [63:0] axi42tl_auto_out_a_bits_data; 
  wire  axi42tl_auto_out_a_bits_corrupt; 
  wire  axi42tl_auto_out_d_ready; 
  wire  axi42tl_auto_out_d_valid; 
  wire [2:0] axi42tl_auto_out_d_bits_opcode; 
  wire [2:0] axi42tl_auto_out_d_bits_size; 
  wire [2:0] axi42tl_auto_out_d_bits_source; 
  wire  axi42tl_auto_out_d_bits_denied; 
  wire [63:0] axi42tl_auto_out_d_bits_data; 
  wire  axi42tl_auto_out_d_bits_corrupt; 
  wire  axi4yank_2_clock; 
  wire  axi4yank_2_reset; 
  wire  axi4yank_2_auto_in_awready; 
  wire  axi4yank_2_auto_in_awvalid; 
  wire  axi4yank_2_auto_in_awid; 
  wire [31:0] axi4yank_2_auto_in_awaddr; 
  wire [7:0] axi4yank_2_auto_in_awlen; 
  wire [2:0] axi4yank_2_auto_in_awsize; 
  wire [16:0] axi4yank_2_auto_in_awuser; 
  wire  axi4yank_2_auto_in_wready; 
  wire  axi4yank_2_auto_in_wvalid; 
  wire [63:0] axi4yank_2_auto_in_wdata; 
  wire [7:0] axi4yank_2_auto_in_wstrb; 
  wire  axi4yank_2_auto_in_wlast; 
  wire  axi4yank_2_auto_in_bready; 
  wire  axi4yank_2_auto_in_bvalid; 
  wire  axi4yank_2_auto_in_bid; 
  wire [1:0] axi4yank_2_auto_in_bresp; 
  wire [16:0] axi4yank_2_auto_in_buser; 
  wire  axi4yank_2_auto_in_arready; 
  wire  axi4yank_2_auto_in_arvalid; 
  wire  axi4yank_2_auto_in_arid; 
  wire [31:0] axi4yank_2_auto_in_araddr; 
  wire [7:0] axi4yank_2_auto_in_arlen; 
  wire [2:0] axi4yank_2_auto_in_arsize; 
  wire [16:0] axi4yank_2_auto_in_aruser; 
  wire  axi4yank_2_auto_in_rready; 
  wire  axi4yank_2_auto_in_rvalid; 
  wire  axi4yank_2_auto_in_rid; 
  wire [63:0] axi4yank_2_auto_in_rdata; 
  wire [1:0] axi4yank_2_auto_in_rresp; 
  wire [16:0] axi4yank_2_auto_in_ruser; 
  wire  axi4yank_2_auto_in_rlast; 
  wire  axi4yank_2_auto_out_awready; 
  wire  axi4yank_2_auto_out_awvalid; 
  wire  axi4yank_2_auto_out_awid; 
  wire [31:0] axi4yank_2_auto_out_awaddr; 
  wire [7:0] axi4yank_2_auto_out_awlen; 
  wire [2:0] axi4yank_2_auto_out_awsize; 
  wire  axi4yank_2_auto_out_wready; 
  wire  axi4yank_2_auto_out_wvalid; 
  wire [63:0] axi4yank_2_auto_out_wdata; 
  wire [7:0] axi4yank_2_auto_out_wstrb; 
  wire  axi4yank_2_auto_out_wlast; 
  wire  axi4yank_2_auto_out_bready; 
  wire  axi4yank_2_auto_out_bvalid; 
  wire  axi4yank_2_auto_out_bid; 
  wire [1:0] axi4yank_2_auto_out_bresp; 
  wire  axi4yank_2_auto_out_arready; 
  wire  axi4yank_2_auto_out_arvalid; 
  wire  axi4yank_2_auto_out_arid; 
  wire [31:0] axi4yank_2_auto_out_araddr; 
  wire [7:0] axi4yank_2_auto_out_arlen; 
  wire [2:0] axi4yank_2_auto_out_arsize; 
  wire  axi4yank_2_auto_out_rready; 
  wire  axi4yank_2_auto_out_rvalid; 
  wire  axi4yank_2_auto_out_rid; 
  wire [63:0] axi4yank_2_auto_out_rdata; 
  wire [1:0] axi4yank_2_auto_out_rresp; 
  wire  axi4yank_2_auto_out_rlast; 
  wire  axi4frag_clock; 
  wire  axi4frag_reset; 
  wire  axi4frag_auto_in_awready; 
  wire  axi4frag_auto_in_awvalid; 
  wire  axi4frag_auto_in_awid; 
  wire [31:0] axi4frag_auto_in_awaddr; 
  wire [7:0] axi4frag_auto_in_awlen; 
  wire [2:0] axi4frag_auto_in_awsize; 
  wire [1:0] axi4frag_auto_in_awburst; 
  wire [15:0] axi4frag_auto_in_awuser; 
  wire  axi4frag_auto_in_wready; 
  wire  axi4frag_auto_in_wvalid; 
  wire [63:0] axi4frag_auto_in_wdata; 
  wire [7:0] axi4frag_auto_in_wstrb; 
  wire  axi4frag_auto_in_wlast; 
  wire  axi4frag_auto_in_bready; 
  wire  axi4frag_auto_in_bvalid; 
  wire  axi4frag_auto_in_bid; 
  wire [1:0] axi4frag_auto_in_bresp; 
  wire [15:0] axi4frag_auto_in_buser; 
  wire  axi4frag_auto_in_arready; 
  wire  axi4frag_auto_in_arvalid; 
  wire  axi4frag_auto_in_arid; 
  wire [31:0] axi4frag_auto_in_araddr; 
  wire [7:0] axi4frag_auto_in_arlen; 
  wire [2:0] axi4frag_auto_in_arsize; 
  wire [1:0] axi4frag_auto_in_arburst; 
  wire [15:0] axi4frag_auto_in_aruser; 
  wire  axi4frag_auto_in_rready; 
  wire  axi4frag_auto_in_rvalid; 
  wire  axi4frag_auto_in_rid; 
  wire [63:0] axi4frag_auto_in_rdata; 
  wire [1:0] axi4frag_auto_in_rresp; 
  wire [15:0] axi4frag_auto_in_ruser; 
  wire  axi4frag_auto_in_rlast; 
  wire  axi4frag_auto_out_awready; 
  wire  axi4frag_auto_out_awvalid; 
  wire  axi4frag_auto_out_awid; 
  wire [31:0] axi4frag_auto_out_awaddr; 
  wire [7:0] axi4frag_auto_out_awlen; 
  wire [2:0] axi4frag_auto_out_awsize; 
  wire [16:0] axi4frag_auto_out_awuser; 
  wire  axi4frag_auto_out_wready; 
  wire  axi4frag_auto_out_wvalid; 
  wire [63:0] axi4frag_auto_out_wdata; 
  wire [7:0] axi4frag_auto_out_wstrb; 
  wire  axi4frag_auto_out_wlast; 
  wire  axi4frag_auto_out_bready; 
  wire  axi4frag_auto_out_bvalid; 
  wire  axi4frag_auto_out_bid; 
  wire [1:0] axi4frag_auto_out_bresp; 
  wire [16:0] axi4frag_auto_out_buser; 
  wire  axi4frag_auto_out_arready; 
  wire  axi4frag_auto_out_arvalid; 
  wire  axi4frag_auto_out_arid; 
  wire [31:0] axi4frag_auto_out_araddr; 
  wire [7:0] axi4frag_auto_out_arlen; 
  wire [2:0] axi4frag_auto_out_arsize; 
  wire [16:0] axi4frag_auto_out_aruser; 
  wire  axi4frag_auto_out_rready; 
  wire  axi4frag_auto_out_rvalid; 
  wire  axi4frag_auto_out_rid; 
  wire [63:0] axi4frag_auto_out_rdata; 
  wire [1:0] axi4frag_auto_out_rresp; 
  wire [16:0] axi4frag_auto_out_ruser; 
  wire  axi4frag_auto_out_rlast; 
  wire  axi4index_2_auto_in_awready; 
  wire  axi4index_2_auto_in_awvalid; 
  wire [16:0] axi4index_2_auto_in_awid; 
  wire [31:0] axi4index_2_auto_in_awaddr; 
  wire [7:0] axi4index_2_auto_in_awlen; 
  wire [2:0] axi4index_2_auto_in_awsize; 
  wire [1:0] axi4index_2_auto_in_awburst; 
  wire  axi4index_2_auto_in_wready; 
  wire  axi4index_2_auto_in_wvalid; 
  wire [63:0] axi4index_2_auto_in_wdata; 
  wire [7:0] axi4index_2_auto_in_wstrb; 
  wire  axi4index_2_auto_in_wlast; 
  wire  axi4index_2_auto_in_bready; 
  wire  axi4index_2_auto_in_bvalid; 
  wire [16:0] axi4index_2_auto_in_bid; 
  wire [1:0] axi4index_2_auto_in_bresp; 
  wire  axi4index_2_auto_in_arready; 
  wire  axi4index_2_auto_in_arvalid; 
  wire [16:0] axi4index_2_auto_in_arid; 
  wire [31:0] axi4index_2_auto_in_araddr; 
  wire [7:0] axi4index_2_auto_in_arlen; 
  wire [2:0] axi4index_2_auto_in_arsize; 
  wire [1:0] axi4index_2_auto_in_arburst; 
  wire  axi4index_2_auto_in_rready; 
  wire  axi4index_2_auto_in_rvalid; 
  wire [16:0] axi4index_2_auto_in_rid; 
  wire [63:0] axi4index_2_auto_in_rdata; 
  wire [1:0] axi4index_2_auto_in_rresp; 
  wire  axi4index_2_auto_in_rlast; 
  wire  axi4index_2_auto_out_awready; 
  wire  axi4index_2_auto_out_awvalid; 
  wire  axi4index_2_auto_out_awid; 
  wire [31:0] axi4index_2_auto_out_awaddr; 
  wire [7:0] axi4index_2_auto_out_awlen; 
  wire [2:0] axi4index_2_auto_out_awsize; 
  wire [1:0] axi4index_2_auto_out_awburst; 
  wire [15:0] axi4index_2_auto_out_awuser; 
  wire  axi4index_2_auto_out_wready; 
  wire  axi4index_2_auto_out_wvalid; 
  wire [63:0] axi4index_2_auto_out_wdata; 
  wire [7:0] axi4index_2_auto_out_wstrb; 
  wire  axi4index_2_auto_out_wlast; 
  wire  axi4index_2_auto_out_bready; 
  wire  axi4index_2_auto_out_bvalid; 
  wire  axi4index_2_auto_out_bid; 
  wire [1:0] axi4index_2_auto_out_bresp; 
  wire [15:0] axi4index_2_auto_out_buser; 
  wire  axi4index_2_auto_out_arready; 
  wire  axi4index_2_auto_out_arvalid; 
  wire  axi4index_2_auto_out_arid; 
  wire [31:0] axi4index_2_auto_out_araddr; 
  wire [7:0] axi4index_2_auto_out_arlen; 
  wire [2:0] axi4index_2_auto_out_arsize; 
  wire [1:0] axi4index_2_auto_out_arburst; 
  wire [15:0] axi4index_2_auto_out_aruser; 
  wire  axi4index_2_auto_out_rready; 
  wire  axi4index_2_auto_out_rvalid; 
  wire  axi4index_2_auto_out_rid; 
  wire [63:0] axi4index_2_auto_out_rdata; 
  wire [1:0] axi4index_2_auto_out_rresp; 
  wire [15:0] axi4index_2_auto_out_ruser; 
  wire  axi4index_2_auto_out_rlast; 
  wire  err_clock; 
  wire  err_reset; 
  wire  err_auto_in_a_ready; 
  wire  err_auto_in_a_valid; 
  wire [2:0] err_auto_in_a_bits_opcode; 
  wire [2:0] err_auto_in_a_bits_param; 
  wire [2:0] err_auto_in_a_bits_size; 
  wire [6:0] err_auto_in_a_bits_source; 
  wire [28:0] err_auto_in_a_bits_address; 
  wire [3:0] err_auto_in_a_bits_mask; 
  wire  err_auto_in_a_bits_corrupt; 
  wire  err_auto_in_c_ready; 
  wire  err_auto_in_c_valid; 
  wire [2:0] err_auto_in_c_bits_opcode; 
  wire [2:0] err_auto_in_c_bits_param; 
  wire [2:0] err_auto_in_c_bits_size; 
  wire [6:0] err_auto_in_c_bits_source; 
  wire [28:0] err_auto_in_c_bits_address; 
  wire  err_auto_in_c_bits_corrupt; 
  wire  err_auto_in_d_ready; 
  wire  err_auto_in_d_valid; 
  wire [2:0] err_auto_in_d_bits_opcode; 
  wire [1:0] err_auto_in_d_bits_param; 
  wire [2:0] err_auto_in_d_bits_size; 
  wire [6:0] err_auto_in_d_bits_source; 
  wire  err_auto_in_d_bits_sink; 
  wire  err_auto_in_d_bits_denied; 
  wire [31:0] err_auto_in_d_bits_data; 
  wire  err_auto_in_d_bits_corrupt; 
  wire  err_auto_in_e_valid; 
  wire  atomics_clock; 
  wire  atomics_reset; 
  wire  atomics_auto_in_a_ready; 
  wire  atomics_auto_in_a_valid; 
  wire [2:0] atomics_auto_in_a_bits_opcode; 
  wire [2:0] atomics_auto_in_a_bits_param; 
  wire [3:0] atomics_auto_in_a_bits_size; 
  wire [6:0] atomics_auto_in_a_bits_source; 
  wire [31:0] atomics_auto_in_a_bits_address; 
  wire [7:0] atomics_auto_in_a_bits_mask; 
  wire [63:0] atomics_auto_in_a_bits_data; 
  wire  atomics_auto_in_c_ready; 
  wire  atomics_auto_in_c_valid; 
  wire [2:0] atomics_auto_in_c_bits_opcode; 
  wire [2:0] atomics_auto_in_c_bits_param; 
  wire [3:0] atomics_auto_in_c_bits_size; 
  wire [6:0] atomics_auto_in_c_bits_source; 
  wire [31:0] atomics_auto_in_c_bits_address; 
  wire  atomics_auto_in_c_bits_corrupt; 
  wire  atomics_auto_in_d_ready; 
  wire  atomics_auto_in_d_valid; 
  wire [2:0] atomics_auto_in_d_bits_opcode; 
  wire [1:0] atomics_auto_in_d_bits_param; 
  wire [3:0] atomics_auto_in_d_bits_size; 
  wire [6:0] atomics_auto_in_d_bits_source; 
  wire  atomics_auto_in_d_bits_sink; 
  wire  atomics_auto_in_d_bits_denied; 
  wire [63:0] atomics_auto_in_d_bits_data; 
  wire  atomics_auto_in_d_bits_corrupt; 
  wire  atomics_auto_in_e_ready; 
  wire  atomics_auto_in_e_valid; 
  wire  atomics_auto_in_e_bits_sink; 
  wire  atomics_auto_out_a_ready; 
  wire  atomics_auto_out_a_valid; 
  wire [2:0] atomics_auto_out_a_bits_opcode; 
  wire [2:0] atomics_auto_out_a_bits_param; 
  wire [3:0] atomics_auto_out_a_bits_size; 
  wire [6:0] atomics_auto_out_a_bits_source; 
  wire [31:0] atomics_auto_out_a_bits_address; 
  wire [7:0] atomics_auto_out_a_bits_mask; 
  wire [63:0] atomics_auto_out_a_bits_data; 
  wire  atomics_auto_out_a_bits_corrupt; 
  wire  atomics_auto_out_c_ready; 
  wire  atomics_auto_out_c_valid; 
  wire [2:0] atomics_auto_out_c_bits_opcode; 
  wire [2:0] atomics_auto_out_c_bits_param; 
  wire [3:0] atomics_auto_out_c_bits_size; 
  wire [6:0] atomics_auto_out_c_bits_source; 
  wire [31:0] atomics_auto_out_c_bits_address; 
  wire  atomics_auto_out_c_bits_corrupt; 
  wire  atomics_auto_out_d_ready; 
  wire  atomics_auto_out_d_valid; 
  wire [2:0] atomics_auto_out_d_bits_opcode; 
  wire [1:0] atomics_auto_out_d_bits_param; 
  wire [3:0] atomics_auto_out_d_bits_size; 
  wire [6:0] atomics_auto_out_d_bits_source; 
  wire  atomics_auto_out_d_bits_sink; 
  wire  atomics_auto_out_d_bits_denied; 
  wire [63:0] atomics_auto_out_d_bits_data; 
  wire  atomics_auto_out_d_bits_corrupt; 
  wire  atomics_auto_out_e_ready; 
  wire  atomics_auto_out_e_valid; 
  wire  atomics_auto_out_e_bits_sink; 
  wire  fixer_1_clock; 
  wire  fixer_1_reset; 
  wire  fixer_1_auto_in_a_ready; 
  wire  fixer_1_auto_in_a_valid; 
  wire [2:0] fixer_1_auto_in_a_bits_opcode; 
  wire [2:0] fixer_1_auto_in_a_bits_param; 
  wire [3:0] fixer_1_auto_in_a_bits_size; 
  wire [6:0] fixer_1_auto_in_a_bits_source; 
  wire [31:0] fixer_1_auto_in_a_bits_address; 
  wire [7:0] fixer_1_auto_in_a_bits_mask; 
  wire [63:0] fixer_1_auto_in_a_bits_data; 
  wire  fixer_1_auto_in_c_ready; 
  wire  fixer_1_auto_in_c_valid; 
  wire [2:0] fixer_1_auto_in_c_bits_opcode; 
  wire [2:0] fixer_1_auto_in_c_bits_param; 
  wire [3:0] fixer_1_auto_in_c_bits_size; 
  wire [6:0] fixer_1_auto_in_c_bits_source; 
  wire [31:0] fixer_1_auto_in_c_bits_address; 
  wire  fixer_1_auto_in_c_bits_corrupt; 
  wire  fixer_1_auto_in_d_ready; 
  wire  fixer_1_auto_in_d_valid; 
  wire [2:0] fixer_1_auto_in_d_bits_opcode; 
  wire [1:0] fixer_1_auto_in_d_bits_param; 
  wire [3:0] fixer_1_auto_in_d_bits_size; 
  wire [6:0] fixer_1_auto_in_d_bits_source; 
  wire  fixer_1_auto_in_d_bits_sink; 
  wire  fixer_1_auto_in_d_bits_denied; 
  wire [63:0] fixer_1_auto_in_d_bits_data; 
  wire  fixer_1_auto_in_d_bits_corrupt; 
  wire  fixer_1_auto_in_e_ready; 
  wire  fixer_1_auto_in_e_valid; 
  wire  fixer_1_auto_in_e_bits_sink; 
  wire  fixer_1_auto_out_a_ready; 
  wire  fixer_1_auto_out_a_valid; 
  wire [2:0] fixer_1_auto_out_a_bits_opcode; 
  wire [2:0] fixer_1_auto_out_a_bits_param; 
  wire [3:0] fixer_1_auto_out_a_bits_size; 
  wire [6:0] fixer_1_auto_out_a_bits_source; 
  wire [31:0] fixer_1_auto_out_a_bits_address; 
  wire [7:0] fixer_1_auto_out_a_bits_mask; 
  wire [63:0] fixer_1_auto_out_a_bits_data; 
  wire  fixer_1_auto_out_c_ready; 
  wire  fixer_1_auto_out_c_valid; 
  wire [2:0] fixer_1_auto_out_c_bits_opcode; 
  wire [2:0] fixer_1_auto_out_c_bits_param; 
  wire [3:0] fixer_1_auto_out_c_bits_size; 
  wire [6:0] fixer_1_auto_out_c_bits_source; 
  wire [31:0] fixer_1_auto_out_c_bits_address; 
  wire  fixer_1_auto_out_c_bits_corrupt; 
  wire  fixer_1_auto_out_d_ready; 
  wire  fixer_1_auto_out_d_valid; 
  wire [2:0] fixer_1_auto_out_d_bits_opcode; 
  wire [1:0] fixer_1_auto_out_d_bits_param; 
  wire [3:0] fixer_1_auto_out_d_bits_size; 
  wire [6:0] fixer_1_auto_out_d_bits_source; 
  wire  fixer_1_auto_out_d_bits_sink; 
  wire  fixer_1_auto_out_d_bits_denied; 
  wire [63:0] fixer_1_auto_out_d_bits_data; 
  wire  fixer_1_auto_out_d_bits_corrupt; 
  wire  fixer_1_auto_out_e_ready; 
  wire  fixer_1_auto_out_e_valid; 
  wire  fixer_1_auto_out_e_bits_sink; 
  wire  hints_clock; 
  wire  hints_reset; 
  wire  hints_auto_in_a_ready; 
  wire  hints_auto_in_a_valid; 
  wire [2:0] hints_auto_in_a_bits_opcode; 
  wire [2:0] hints_auto_in_a_bits_param; 
  wire [3:0] hints_auto_in_a_bits_size; 
  wire [5:0] hints_auto_in_a_bits_source; 
  wire [31:0] hints_auto_in_a_bits_address; 
  wire [7:0] hints_auto_in_a_bits_mask; 
  wire [63:0] hints_auto_in_a_bits_data; 
  wire  hints_auto_in_c_ready; 
  wire  hints_auto_in_c_valid; 
  wire [2:0] hints_auto_in_c_bits_opcode; 
  wire [2:0] hints_auto_in_c_bits_param; 
  wire [3:0] hints_auto_in_c_bits_size; 
  wire [5:0] hints_auto_in_c_bits_source; 
  wire [31:0] hints_auto_in_c_bits_address; 
  wire  hints_auto_in_c_bits_corrupt; 
  wire  hints_auto_in_d_ready; 
  wire  hints_auto_in_d_valid; 
  wire [2:0] hints_auto_in_d_bits_opcode; 
  wire [1:0] hints_auto_in_d_bits_param; 
  wire [3:0] hints_auto_in_d_bits_size; 
  wire [5:0] hints_auto_in_d_bits_source; 
  wire  hints_auto_in_d_bits_sink; 
  wire  hints_auto_in_d_bits_denied; 
  wire [63:0] hints_auto_in_d_bits_data; 
  wire  hints_auto_in_d_bits_corrupt; 
  wire  hints_auto_in_e_ready; 
  wire  hints_auto_in_e_valid; 
  wire  hints_auto_in_e_bits_sink; 
  wire  hints_auto_out_a_ready; 
  wire  hints_auto_out_a_valid; 
  wire [2:0] hints_auto_out_a_bits_opcode; 
  wire [2:0] hints_auto_out_a_bits_param; 
  wire [3:0] hints_auto_out_a_bits_size; 
  wire [6:0] hints_auto_out_a_bits_source; 
  wire [31:0] hints_auto_out_a_bits_address; 
  wire [7:0] hints_auto_out_a_bits_mask; 
  wire [63:0] hints_auto_out_a_bits_data; 
  wire  hints_auto_out_c_ready; 
  wire  hints_auto_out_c_valid; 
  wire [2:0] hints_auto_out_c_bits_opcode; 
  wire [2:0] hints_auto_out_c_bits_param; 
  wire [3:0] hints_auto_out_c_bits_size; 
  wire [6:0] hints_auto_out_c_bits_source; 
  wire [31:0] hints_auto_out_c_bits_address; 
  wire  hints_auto_out_c_bits_corrupt; 
  wire  hints_auto_out_d_ready; 
  wire  hints_auto_out_d_valid; 
  wire [2:0] hints_auto_out_d_bits_opcode; 
  wire [1:0] hints_auto_out_d_bits_param; 
  wire [3:0] hints_auto_out_d_bits_size; 
  wire [6:0] hints_auto_out_d_bits_source; 
  wire  hints_auto_out_d_bits_sink; 
  wire  hints_auto_out_d_bits_denied; 
  wire [63:0] hints_auto_out_d_bits_data; 
  wire  hints_auto_out_d_bits_corrupt; 
  wire  hints_auto_out_e_ready; 
  wire  hints_auto_out_e_valid; 
  wire  hints_auto_out_e_bits_sink; 
  wire  widget_1_clock; 
  wire  widget_1_reset; 
  wire  widget_1_auto_in_a_ready; 
  wire  widget_1_auto_in_a_valid; 
  wire [2:0] widget_1_auto_in_a_bits_opcode; 
  wire [2:0] widget_1_auto_in_a_bits_param; 
  wire [3:0] widget_1_auto_in_a_bits_size; 
  wire [5:0] widget_1_auto_in_a_bits_source; 
  wire [31:0] widget_1_auto_in_a_bits_address; 
  wire [3:0] widget_1_auto_in_a_bits_mask; 
  wire [31:0] widget_1_auto_in_a_bits_data; 
  wire  widget_1_auto_in_c_ready; 
  wire  widget_1_auto_in_c_valid; 
  wire [2:0] widget_1_auto_in_c_bits_opcode; 
  wire [2:0] widget_1_auto_in_c_bits_param; 
  wire [3:0] widget_1_auto_in_c_bits_size; 
  wire [5:0] widget_1_auto_in_c_bits_source; 
  wire [31:0] widget_1_auto_in_c_bits_address; 
  wire  widget_1_auto_in_c_bits_corrupt; 
  wire  widget_1_auto_in_d_ready; 
  wire  widget_1_auto_in_d_valid; 
  wire [2:0] widget_1_auto_in_d_bits_opcode; 
  wire [1:0] widget_1_auto_in_d_bits_param; 
  wire [3:0] widget_1_auto_in_d_bits_size; 
  wire [5:0] widget_1_auto_in_d_bits_source; 
  wire  widget_1_auto_in_d_bits_sink; 
  wire  widget_1_auto_in_d_bits_denied; 
  wire [31:0] widget_1_auto_in_d_bits_data; 
  wire  widget_1_auto_in_d_bits_corrupt; 
  wire  widget_1_auto_in_e_ready; 
  wire  widget_1_auto_in_e_valid; 
  wire  widget_1_auto_in_e_bits_sink; 
  wire  widget_1_auto_out_a_ready; 
  wire  widget_1_auto_out_a_valid; 
  wire [2:0] widget_1_auto_out_a_bits_opcode; 
  wire [2:0] widget_1_auto_out_a_bits_param; 
  wire [3:0] widget_1_auto_out_a_bits_size; 
  wire [5:0] widget_1_auto_out_a_bits_source; 
  wire [31:0] widget_1_auto_out_a_bits_address; 
  wire [7:0] widget_1_auto_out_a_bits_mask; 
  wire [63:0] widget_1_auto_out_a_bits_data; 
  wire  widget_1_auto_out_c_ready; 
  wire  widget_1_auto_out_c_valid; 
  wire [2:0] widget_1_auto_out_c_bits_opcode; 
  wire [2:0] widget_1_auto_out_c_bits_param; 
  wire [3:0] widget_1_auto_out_c_bits_size; 
  wire [5:0] widget_1_auto_out_c_bits_source; 
  wire [31:0] widget_1_auto_out_c_bits_address; 
  wire  widget_1_auto_out_c_bits_corrupt; 
  wire  widget_1_auto_out_d_ready; 
  wire  widget_1_auto_out_d_valid; 
  wire [2:0] widget_1_auto_out_d_bits_opcode; 
  wire [1:0] widget_1_auto_out_d_bits_param; 
  wire [3:0] widget_1_auto_out_d_bits_size; 
  wire [5:0] widget_1_auto_out_d_bits_source; 
  wire  widget_1_auto_out_d_bits_sink; 
  wire  widget_1_auto_out_d_bits_denied; 
  wire [63:0] widget_1_auto_out_d_bits_data; 
  wire  widget_1_auto_out_d_bits_corrupt; 
  wire  widget_1_auto_out_e_ready; 
  wire  widget_1_auto_out_e_valid; 
  wire  widget_1_auto_out_e_bits_sink; 
  wire  widget_2_clock; 
  wire  widget_2_reset; 
  wire  widget_2_auto_in_a_ready; 
  wire  widget_2_auto_in_a_valid; 
  wire [2:0] widget_2_auto_in_a_bits_opcode; 
  wire [2:0] widget_2_auto_in_a_bits_param; 
  wire [2:0] widget_2_auto_in_a_bits_size; 
  wire [6:0] widget_2_auto_in_a_bits_source; 
  wire [28:0] widget_2_auto_in_a_bits_address; 
  wire [7:0] widget_2_auto_in_a_bits_mask; 
  wire  widget_2_auto_in_a_bits_corrupt; 
  wire  widget_2_auto_in_c_ready; 
  wire  widget_2_auto_in_c_valid; 
  wire [2:0] widget_2_auto_in_c_bits_opcode; 
  wire [2:0] widget_2_auto_in_c_bits_param; 
  wire [2:0] widget_2_auto_in_c_bits_size; 
  wire [6:0] widget_2_auto_in_c_bits_source; 
  wire [28:0] widget_2_auto_in_c_bits_address; 
  wire  widget_2_auto_in_c_bits_corrupt; 
  wire  widget_2_auto_in_d_ready; 
  wire  widget_2_auto_in_d_valid; 
  wire [2:0] widget_2_auto_in_d_bits_opcode; 
  wire [1:0] widget_2_auto_in_d_bits_param; 
  wire [2:0] widget_2_auto_in_d_bits_size; 
  wire [6:0] widget_2_auto_in_d_bits_source; 
  wire  widget_2_auto_in_d_bits_sink; 
  wire  widget_2_auto_in_d_bits_denied; 
  wire [63:0] widget_2_auto_in_d_bits_data; 
  wire  widget_2_auto_in_d_bits_corrupt; 
  wire  widget_2_auto_in_e_valid; 
  wire  widget_2_auto_out_a_ready; 
  wire  widget_2_auto_out_a_valid; 
  wire [2:0] widget_2_auto_out_a_bits_opcode; 
  wire [2:0] widget_2_auto_out_a_bits_param; 
  wire [2:0] widget_2_auto_out_a_bits_size; 
  wire [6:0] widget_2_auto_out_a_bits_source; 
  wire [28:0] widget_2_auto_out_a_bits_address; 
  wire [3:0] widget_2_auto_out_a_bits_mask; 
  wire  widget_2_auto_out_a_bits_corrupt; 
  wire  widget_2_auto_out_c_ready; 
  wire  widget_2_auto_out_c_valid; 
  wire [2:0] widget_2_auto_out_c_bits_opcode; 
  wire [2:0] widget_2_auto_out_c_bits_param; 
  wire [2:0] widget_2_auto_out_c_bits_size; 
  wire [6:0] widget_2_auto_out_c_bits_source; 
  wire [28:0] widget_2_auto_out_c_bits_address; 
  wire  widget_2_auto_out_c_bits_corrupt; 
  wire  widget_2_auto_out_d_ready; 
  wire  widget_2_auto_out_d_valid; 
  wire [2:0] widget_2_auto_out_d_bits_opcode; 
  wire [1:0] widget_2_auto_out_d_bits_param; 
  wire [2:0] widget_2_auto_out_d_bits_size; 
  wire [6:0] widget_2_auto_out_d_bits_source; 
  wire  widget_2_auto_out_d_bits_sink; 
  wire  widget_2_auto_out_d_bits_denied; 
  wire [31:0] widget_2_auto_out_d_bits_data; 
  wire  widget_2_auto_out_d_bits_corrupt; 
  wire  widget_2_auto_out_e_valid; 
  dual_TLXbar xbar ( 
    .clock(xbar_clock),
    .reset(xbar_reset),
    .auto_in_a_ready(xbar_auto_in_a_ready),
    .auto_in_a_valid(xbar_auto_in_a_valid),
    .auto_in_a_bits_opcode(xbar_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(xbar_auto_in_a_bits_param),
    .auto_in_a_bits_size(xbar_auto_in_a_bits_size),
    .auto_in_a_bits_source(xbar_auto_in_a_bits_source),
    .auto_in_a_bits_address(xbar_auto_in_a_bits_address),
    .auto_in_a_bits_mask(xbar_auto_in_a_bits_mask),
    .auto_in_a_bits_data(xbar_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(xbar_auto_in_a_bits_corrupt),
    .auto_in_c_ready(xbar_auto_in_c_ready),
    .auto_in_c_valid(xbar_auto_in_c_valid),
    .auto_in_c_bits_opcode(xbar_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(xbar_auto_in_c_bits_param),
    .auto_in_c_bits_size(xbar_auto_in_c_bits_size),
    .auto_in_c_bits_source(xbar_auto_in_c_bits_source),
    .auto_in_c_bits_address(xbar_auto_in_c_bits_address),
    .auto_in_c_bits_corrupt(xbar_auto_in_c_bits_corrupt),
    .auto_in_d_ready(xbar_auto_in_d_ready),
    .auto_in_d_valid(xbar_auto_in_d_valid),
    .auto_in_d_bits_opcode(xbar_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(xbar_auto_in_d_bits_param),
    .auto_in_d_bits_size(xbar_auto_in_d_bits_size),
    .auto_in_d_bits_source(xbar_auto_in_d_bits_source),
    .auto_in_d_bits_sink(xbar_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(xbar_auto_in_d_bits_denied),
    .auto_in_d_bits_data(xbar_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(xbar_auto_in_d_bits_corrupt),
    .auto_in_e_ready(xbar_auto_in_e_ready),
    .auto_in_e_valid(xbar_auto_in_e_valid),
    .auto_in_e_bits_sink(xbar_auto_in_e_bits_sink),
    .auto_out_2_a_ready(xbar_auto_out_2_a_ready),
    .auto_out_2_a_valid(xbar_auto_out_2_a_valid),
    .auto_out_2_a_bits_opcode(xbar_auto_out_2_a_bits_opcode),
    .auto_out_2_a_bits_param(xbar_auto_out_2_a_bits_param),
    .auto_out_2_a_bits_size(xbar_auto_out_2_a_bits_size),
    .auto_out_2_a_bits_source(xbar_auto_out_2_a_bits_source),
    .auto_out_2_a_bits_address(xbar_auto_out_2_a_bits_address),
    .auto_out_2_a_bits_mask(xbar_auto_out_2_a_bits_mask),
    .auto_out_2_a_bits_corrupt(xbar_auto_out_2_a_bits_corrupt),
    .auto_out_2_c_ready(xbar_auto_out_2_c_ready),
    .auto_out_2_c_valid(xbar_auto_out_2_c_valid),
    .auto_out_2_c_bits_opcode(xbar_auto_out_2_c_bits_opcode),
    .auto_out_2_c_bits_param(xbar_auto_out_2_c_bits_param),
    .auto_out_2_c_bits_size(xbar_auto_out_2_c_bits_size),
    .auto_out_2_c_bits_source(xbar_auto_out_2_c_bits_source),
    .auto_out_2_c_bits_address(xbar_auto_out_2_c_bits_address),
    .auto_out_2_c_bits_corrupt(xbar_auto_out_2_c_bits_corrupt),
    .auto_out_2_d_ready(xbar_auto_out_2_d_ready),
    .auto_out_2_d_valid(xbar_auto_out_2_d_valid),
    .auto_out_2_d_bits_opcode(xbar_auto_out_2_d_bits_opcode),
    .auto_out_2_d_bits_param(xbar_auto_out_2_d_bits_param),
    .auto_out_2_d_bits_size(xbar_auto_out_2_d_bits_size),
    .auto_out_2_d_bits_source(xbar_auto_out_2_d_bits_source),
    .auto_out_2_d_bits_sink(xbar_auto_out_2_d_bits_sink),
    .auto_out_2_d_bits_denied(xbar_auto_out_2_d_bits_denied),
    .auto_out_2_d_bits_data(xbar_auto_out_2_d_bits_data),
    .auto_out_2_d_bits_corrupt(xbar_auto_out_2_d_bits_corrupt),
    .auto_out_2_e_valid(xbar_auto_out_2_e_valid),
    .auto_out_1_a_ready(xbar_auto_out_1_a_ready),
    .auto_out_1_a_valid(xbar_auto_out_1_a_valid),
    .auto_out_1_a_bits_opcode(xbar_auto_out_1_a_bits_opcode),
    .auto_out_1_a_bits_param(xbar_auto_out_1_a_bits_param),
    .auto_out_1_a_bits_size(xbar_auto_out_1_a_bits_size),
    .auto_out_1_a_bits_source(xbar_auto_out_1_a_bits_source),
    .auto_out_1_a_bits_address(xbar_auto_out_1_a_bits_address),
    .auto_out_1_a_bits_mask(xbar_auto_out_1_a_bits_mask),
    .auto_out_1_a_bits_data(xbar_auto_out_1_a_bits_data),
    .auto_out_1_a_bits_corrupt(xbar_auto_out_1_a_bits_corrupt),
    .auto_out_1_d_ready(xbar_auto_out_1_d_ready),
    .auto_out_1_d_valid(xbar_auto_out_1_d_valid),
    .auto_out_1_d_bits_opcode(xbar_auto_out_1_d_bits_opcode),
    .auto_out_1_d_bits_size(xbar_auto_out_1_d_bits_size),
    .auto_out_1_d_bits_source(xbar_auto_out_1_d_bits_source),
    .auto_out_1_d_bits_denied(xbar_auto_out_1_d_bits_denied),
    .auto_out_1_d_bits_data(xbar_auto_out_1_d_bits_data),
    .auto_out_1_d_bits_corrupt(xbar_auto_out_1_d_bits_corrupt),
    .auto_out_0_a_ready(xbar_auto_out_0_a_ready),
    .auto_out_0_a_valid(xbar_auto_out_0_a_valid),
    .auto_out_0_a_bits_opcode(xbar_auto_out_0_a_bits_opcode),
    .auto_out_0_a_bits_param(xbar_auto_out_0_a_bits_param),
    .auto_out_0_a_bits_size(xbar_auto_out_0_a_bits_size),
    .auto_out_0_a_bits_source(xbar_auto_out_0_a_bits_source),
    .auto_out_0_a_bits_address(xbar_auto_out_0_a_bits_address),
    .auto_out_0_a_bits_mask(xbar_auto_out_0_a_bits_mask),
    .auto_out_0_a_bits_data(xbar_auto_out_0_a_bits_data),
    .auto_out_0_a_bits_corrupt(xbar_auto_out_0_a_bits_corrupt),
    .auto_out_0_d_ready(xbar_auto_out_0_d_ready),
    .auto_out_0_d_valid(xbar_auto_out_0_d_valid),
    .auto_out_0_d_bits_opcode(xbar_auto_out_0_d_bits_opcode),
    .auto_out_0_d_bits_size(xbar_auto_out_0_d_bits_size),
    .auto_out_0_d_bits_source(xbar_auto_out_0_d_bits_source),
    .auto_out_0_d_bits_denied(xbar_auto_out_0_d_bits_denied),
    .auto_out_0_d_bits_data(xbar_auto_out_0_d_bits_data),
    .auto_out_0_d_bits_corrupt(xbar_auto_out_0_d_bits_corrupt)
  );
  dual_TLXbar_1 xbar_1 ( 
    .clock(xbar_1_clock),
    .reset(xbar_1_reset),
    .auto_in_a_ready(xbar_1_auto_in_a_ready),
    .auto_in_a_valid(xbar_1_auto_in_a_valid),
    .auto_in_a_bits_opcode(xbar_1_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(xbar_1_auto_in_a_bits_param),
    .auto_in_a_bits_size(xbar_1_auto_in_a_bits_size),
    .auto_in_a_bits_source(xbar_1_auto_in_a_bits_source),
    .auto_in_a_bits_address(xbar_1_auto_in_a_bits_address),
    .auto_in_a_bits_mask(xbar_1_auto_in_a_bits_mask),
    .auto_in_a_bits_data(xbar_1_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(xbar_1_auto_in_a_bits_corrupt),
    .auto_in_d_ready(xbar_1_auto_in_d_ready),
    .auto_in_d_valid(xbar_1_auto_in_d_valid),
    .auto_in_d_bits_opcode(xbar_1_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(xbar_1_auto_in_d_bits_param),
    .auto_in_d_bits_size(xbar_1_auto_in_d_bits_size),
    .auto_in_d_bits_source(xbar_1_auto_in_d_bits_source),
    .auto_in_d_bits_sink(xbar_1_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(xbar_1_auto_in_d_bits_denied),
    .auto_in_d_bits_data(xbar_1_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(xbar_1_auto_in_d_bits_corrupt),
    .auto_out_1_a_ready(xbar_1_auto_out_1_a_ready),
    .auto_out_1_a_valid(xbar_1_auto_out_1_a_valid),
    .auto_out_1_a_bits_opcode(xbar_1_auto_out_1_a_bits_opcode),
    .auto_out_1_a_bits_param(xbar_1_auto_out_1_a_bits_param),
    .auto_out_1_a_bits_size(xbar_1_auto_out_1_a_bits_size),
    .auto_out_1_a_bits_source(xbar_1_auto_out_1_a_bits_source),
    .auto_out_1_a_bits_address(xbar_1_auto_out_1_a_bits_address),
    .auto_out_1_a_bits_mask(xbar_1_auto_out_1_a_bits_mask),
    .auto_out_1_a_bits_corrupt(xbar_1_auto_out_1_a_bits_corrupt),
    .auto_out_1_d_ready(xbar_1_auto_out_1_d_ready),
    .auto_out_1_d_valid(xbar_1_auto_out_1_d_valid),
    .auto_out_1_d_bits_opcode(xbar_1_auto_out_1_d_bits_opcode),
    .auto_out_1_d_bits_param(xbar_1_auto_out_1_d_bits_param),
    .auto_out_1_d_bits_size(xbar_1_auto_out_1_d_bits_size),
    .auto_out_1_d_bits_source(xbar_1_auto_out_1_d_bits_source),
    .auto_out_1_d_bits_sink(xbar_1_auto_out_1_d_bits_sink),
    .auto_out_1_d_bits_denied(xbar_1_auto_out_1_d_bits_denied),
    .auto_out_1_d_bits_data(xbar_1_auto_out_1_d_bits_data),
    .auto_out_1_d_bits_corrupt(xbar_1_auto_out_1_d_bits_corrupt),
    .auto_out_0_a_ready(xbar_1_auto_out_0_a_ready),
    .auto_out_0_a_valid(xbar_1_auto_out_0_a_valid),
    .auto_out_0_a_bits_opcode(xbar_1_auto_out_0_a_bits_opcode),
    .auto_out_0_a_bits_param(xbar_1_auto_out_0_a_bits_param),
    .auto_out_0_a_bits_size(xbar_1_auto_out_0_a_bits_size),
    .auto_out_0_a_bits_source(xbar_1_auto_out_0_a_bits_source),
    .auto_out_0_a_bits_address(xbar_1_auto_out_0_a_bits_address),
    .auto_out_0_a_bits_mask(xbar_1_auto_out_0_a_bits_mask),
    .auto_out_0_a_bits_data(xbar_1_auto_out_0_a_bits_data),
    .auto_out_0_a_bits_corrupt(xbar_1_auto_out_0_a_bits_corrupt),
    .auto_out_0_d_ready(xbar_1_auto_out_0_d_ready),
    .auto_out_0_d_valid(xbar_1_auto_out_0_d_valid),
    .auto_out_0_d_bits_opcode(xbar_1_auto_out_0_d_bits_opcode),
    .auto_out_0_d_bits_param(xbar_1_auto_out_0_d_bits_param),
    .auto_out_0_d_bits_size(xbar_1_auto_out_0_d_bits_size),
    .auto_out_0_d_bits_source(xbar_1_auto_out_0_d_bits_source),
    .auto_out_0_d_bits_sink(xbar_1_auto_out_0_d_bits_sink),
    .auto_out_0_d_bits_denied(xbar_1_auto_out_0_d_bits_denied),
    .auto_out_0_d_bits_data(xbar_1_auto_out_0_d_bits_data),
    .auto_out_0_d_bits_corrupt(xbar_1_auto_out_0_d_bits_corrupt)
  );
  dual_TLError ferr ( 
    .clock(ferr_clock),
    .reset(ferr_reset),
    .auto_in_a_ready(ferr_auto_in_a_ready),
    .auto_in_a_valid(ferr_auto_in_a_valid),
    .auto_in_a_bits_opcode(ferr_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(ferr_auto_in_a_bits_param),
    .auto_in_a_bits_size(ferr_auto_in_a_bits_size),
    .auto_in_a_bits_source(ferr_auto_in_a_bits_source),
    .auto_in_a_bits_address(ferr_auto_in_a_bits_address),
    .auto_in_a_bits_mask(ferr_auto_in_a_bits_mask),
    .auto_in_a_bits_corrupt(ferr_auto_in_a_bits_corrupt),
    .auto_in_d_ready(ferr_auto_in_d_ready),
    .auto_in_d_valid(ferr_auto_in_d_valid),
    .auto_in_d_bits_opcode(ferr_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(ferr_auto_in_d_bits_param),
    .auto_in_d_bits_size(ferr_auto_in_d_bits_size),
    .auto_in_d_bits_source(ferr_auto_in_d_bits_source),
    .auto_in_d_bits_sink(ferr_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(ferr_auto_in_d_bits_denied),
    .auto_in_d_bits_data(ferr_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(ferr_auto_in_d_bits_corrupt)
  );
  dual_ChipLink chiplink ( 
    .clock(chiplink_clock),
    .reset(chiplink_reset),
    .auto_mbypass_out_a_ready(chiplink_auto_mbypass_out_a_ready),
    .auto_mbypass_out_a_valid(chiplink_auto_mbypass_out_a_valid),
    .auto_mbypass_out_a_bits_opcode(chiplink_auto_mbypass_out_a_bits_opcode),
    .auto_mbypass_out_a_bits_param(chiplink_auto_mbypass_out_a_bits_param),
    .auto_mbypass_out_a_bits_size(chiplink_auto_mbypass_out_a_bits_size),
    .auto_mbypass_out_a_bits_source(chiplink_auto_mbypass_out_a_bits_source),
    .auto_mbypass_out_a_bits_address(chiplink_auto_mbypass_out_a_bits_address),
    .auto_mbypass_out_a_bits_mask(chiplink_auto_mbypass_out_a_bits_mask),
    .auto_mbypass_out_a_bits_data(chiplink_auto_mbypass_out_a_bits_data),
    .auto_mbypass_out_c_ready(chiplink_auto_mbypass_out_c_ready),
    .auto_mbypass_out_c_valid(chiplink_auto_mbypass_out_c_valid),
    .auto_mbypass_out_c_bits_opcode(chiplink_auto_mbypass_out_c_bits_opcode),
    .auto_mbypass_out_c_bits_param(chiplink_auto_mbypass_out_c_bits_param),
    .auto_mbypass_out_c_bits_size(chiplink_auto_mbypass_out_c_bits_size),
    .auto_mbypass_out_c_bits_source(chiplink_auto_mbypass_out_c_bits_source),
    .auto_mbypass_out_c_bits_address(chiplink_auto_mbypass_out_c_bits_address),
    .auto_mbypass_out_c_bits_corrupt(chiplink_auto_mbypass_out_c_bits_corrupt),
    .auto_mbypass_out_d_ready(chiplink_auto_mbypass_out_d_ready),
    .auto_mbypass_out_d_valid(chiplink_auto_mbypass_out_d_valid),
    .auto_mbypass_out_d_bits_opcode(chiplink_auto_mbypass_out_d_bits_opcode),
    .auto_mbypass_out_d_bits_param(chiplink_auto_mbypass_out_d_bits_param),
    .auto_mbypass_out_d_bits_size(chiplink_auto_mbypass_out_d_bits_size),
    .auto_mbypass_out_d_bits_source(chiplink_auto_mbypass_out_d_bits_source),
    .auto_mbypass_out_d_bits_sink(chiplink_auto_mbypass_out_d_bits_sink),
    .auto_mbypass_out_d_bits_denied(chiplink_auto_mbypass_out_d_bits_denied),
    .auto_mbypass_out_d_bits_data(chiplink_auto_mbypass_out_d_bits_data),
    .auto_mbypass_out_d_bits_corrupt(chiplink_auto_mbypass_out_d_bits_corrupt),
    .auto_mbypass_out_e_ready(chiplink_auto_mbypass_out_e_ready),
    .auto_mbypass_out_e_valid(chiplink_auto_mbypass_out_e_valid),
    .auto_mbypass_out_e_bits_sink(chiplink_auto_mbypass_out_e_bits_sink),
    .auto_sbypass_node_in_in_a_ready(chiplink_auto_sbypass_node_in_in_a_ready),
    .auto_sbypass_node_in_in_a_valid(chiplink_auto_sbypass_node_in_in_a_valid),
    .auto_sbypass_node_in_in_a_bits_opcode(chiplink_auto_sbypass_node_in_in_a_bits_opcode),
    .auto_sbypass_node_in_in_a_bits_param(chiplink_auto_sbypass_node_in_in_a_bits_param),
    .auto_sbypass_node_in_in_a_bits_size(chiplink_auto_sbypass_node_in_in_a_bits_size),
    .auto_sbypass_node_in_in_a_bits_source(chiplink_auto_sbypass_node_in_in_a_bits_source),
    .auto_sbypass_node_in_in_a_bits_address(chiplink_auto_sbypass_node_in_in_a_bits_address),
    .auto_sbypass_node_in_in_a_bits_mask(chiplink_auto_sbypass_node_in_in_a_bits_mask),
    .auto_sbypass_node_in_in_a_bits_data(chiplink_auto_sbypass_node_in_in_a_bits_data),
    .auto_sbypass_node_in_in_a_bits_corrupt(chiplink_auto_sbypass_node_in_in_a_bits_corrupt),
    .auto_sbypass_node_in_in_d_ready(chiplink_auto_sbypass_node_in_in_d_ready),
    .auto_sbypass_node_in_in_d_valid(chiplink_auto_sbypass_node_in_in_d_valid),
    .auto_sbypass_node_in_in_d_bits_opcode(chiplink_auto_sbypass_node_in_in_d_bits_opcode),
    .auto_sbypass_node_in_in_d_bits_param(chiplink_auto_sbypass_node_in_in_d_bits_param),
    .auto_sbypass_node_in_in_d_bits_size(chiplink_auto_sbypass_node_in_in_d_bits_size),
    .auto_sbypass_node_in_in_d_bits_source(chiplink_auto_sbypass_node_in_in_d_bits_source),
    .auto_sbypass_node_in_in_d_bits_sink(chiplink_auto_sbypass_node_in_in_d_bits_sink),
    .auto_sbypass_node_in_in_d_bits_denied(chiplink_auto_sbypass_node_in_in_d_bits_denied),
    .auto_sbypass_node_in_in_d_bits_data(chiplink_auto_sbypass_node_in_in_d_bits_data),
    .auto_sbypass_node_in_in_d_bits_corrupt(chiplink_auto_sbypass_node_in_in_d_bits_corrupt),
    .auto_io_out_c2b_clk(chiplink_auto_io_out_c2b_clk),
    .auto_io_out_c2b_rst(chiplink_auto_io_out_c2b_rst),
    .auto_io_out_c2b_send(chiplink_auto_io_out_c2b_send),
    .auto_io_out_c2b_data(chiplink_auto_io_out_c2b_data),
    .auto_io_out_b2c_clk(chiplink_auto_io_out_b2c_clk),
    .auto_io_out_b2c_rst(chiplink_auto_io_out_b2c_rst),
    .auto_io_out_b2c_send(chiplink_auto_io_out_b2c_send),
    .auto_io_out_b2c_data(chiplink_auto_io_out_b2c_data)
  );
  dual_AXI4UserYanker axi4yank ( 
    .clock(axi4yank_clock),
    .reset(axi4yank_reset),
    .auto_in_awready(axi4yank_auto_in_awready),
    .auto_in_awvalid(axi4yank_auto_in_awvalid),
    .auto_in_awid(axi4yank_auto_in_awid),
    .auto_in_awaddr(axi4yank_auto_in_awaddr),
    .auto_in_awlen(axi4yank_auto_in_awlen),
    .auto_in_awsize(axi4yank_auto_in_awsize),
    .auto_in_awburst(axi4yank_auto_in_awburst),
    .auto_in_awlock(axi4yank_auto_in_awlock),
    .auto_in_awcache(axi4yank_auto_in_awcache),
    .auto_in_awprot(axi4yank_auto_in_awprot),
    .auto_in_awqos(axi4yank_auto_in_awqos),
    .auto_in_awuser(axi4yank_auto_in_awuser),
    .auto_in_awinstret(axi4yank_auto_in_awinstret),
    .auto_in_wready(axi4yank_auto_in_wready),
    .auto_in_wvalid(axi4yank_auto_in_wvalid),
    .auto_in_wdata(axi4yank_auto_in_wdata),
    .auto_in_wstrb(axi4yank_auto_in_wstrb),
    .auto_in_wlast(axi4yank_auto_in_wlast),
    .auto_in_bready(axi4yank_auto_in_bready),
    .auto_in_bvalid(axi4yank_auto_in_bvalid),
    .auto_in_bid(axi4yank_auto_in_bid),
    .auto_in_bresp(axi4yank_auto_in_bresp),
    .auto_in_buser(axi4yank_auto_in_buser),
    .auto_in_arready(axi4yank_auto_in_arready),
    .auto_in_arvalid(axi4yank_auto_in_arvalid),
    .auto_in_arid(axi4yank_auto_in_arid),
    .auto_in_araddr(axi4yank_auto_in_araddr),
    .auto_in_arlen(axi4yank_auto_in_arlen),
    .auto_in_arsize(axi4yank_auto_in_arsize),
    .auto_in_arburst(axi4yank_auto_in_arburst),
    .auto_in_arlock(axi4yank_auto_in_arlock),
    .auto_in_arcache(axi4yank_auto_in_arcache),
    .auto_in_arprot(axi4yank_auto_in_arprot),
    .auto_in_arqos(axi4yank_auto_in_arqos),
    .auto_in_aruser(axi4yank_auto_in_aruser),
    .auto_in_arinstret(axi4yank_auto_in_arinstret),
    .auto_in_rready(axi4yank_auto_in_rready),
    .auto_in_rvalid(axi4yank_auto_in_rvalid),
    .auto_in_rid(axi4yank_auto_in_rid),
    .auto_in_rdata(axi4yank_auto_in_rdata),
    .auto_in_rresp(axi4yank_auto_in_rresp),
    .auto_in_ruser(axi4yank_auto_in_ruser),
    .auto_in_rlast(axi4yank_auto_in_rlast),
    .auto_out_awready(axi4yank_auto_out_awready),
    .auto_out_awvalid(axi4yank_auto_out_awvalid),
    .auto_out_awid(axi4yank_auto_out_awid),
    .auto_out_awaddr(axi4yank_auto_out_awaddr),
    .auto_out_awlen(axi4yank_auto_out_awlen),
    .auto_out_awsize(axi4yank_auto_out_awsize),
    .auto_out_awburst(axi4yank_auto_out_awburst),
    .auto_out_awlock(axi4yank_auto_out_awlock),
    .auto_out_awcache(axi4yank_auto_out_awcache),
    .auto_out_awprot(axi4yank_auto_out_awprot),
    .auto_out_awqos(axi4yank_auto_out_awqos),
    .auto_out_awinstret(axi4yank_auto_out_awinstret),
    .auto_out_wready(axi4yank_auto_out_wready),
    .auto_out_wvalid(axi4yank_auto_out_wvalid),
    .auto_out_wdata(axi4yank_auto_out_wdata),
    .auto_out_wstrb(axi4yank_auto_out_wstrb),
    .auto_out_wlast(axi4yank_auto_out_wlast),
    .auto_out_bready(axi4yank_auto_out_bready),
    .auto_out_bvalid(axi4yank_auto_out_bvalid),
    .auto_out_bid(axi4yank_auto_out_bid),
    .auto_out_bresp(axi4yank_auto_out_bresp),
    .auto_out_arready(axi4yank_auto_out_arready),
    .auto_out_arvalid(axi4yank_auto_out_arvalid),
    .auto_out_arid(axi4yank_auto_out_arid),
    .auto_out_araddr(axi4yank_auto_out_araddr),
    .auto_out_arlen(axi4yank_auto_out_arlen),
    .auto_out_arsize(axi4yank_auto_out_arsize),
    .auto_out_arburst(axi4yank_auto_out_arburst),
    .auto_out_arlock(axi4yank_auto_out_arlock),
    .auto_out_arcache(axi4yank_auto_out_arcache),
    .auto_out_arprot(axi4yank_auto_out_arprot),
    .auto_out_arqos(axi4yank_auto_out_arqos),
    .auto_out_arinstret(axi4yank_auto_out_arinstret),
    .auto_out_rready(axi4yank_auto_out_rready),
    .auto_out_rvalid(axi4yank_auto_out_rvalid),
    .auto_out_rid(axi4yank_auto_out_rid),
    .auto_out_rdata(axi4yank_auto_out_rdata),
    .auto_out_rresp(axi4yank_auto_out_rresp),
    .auto_out_rlast(axi4yank_auto_out_rlast)
  );
  dual_AXI4IdIndexer axi4index ( 
    .auto_in_awready(axi4index_auto_in_awready),
    .auto_in_awvalid(axi4index_auto_in_awvalid),
    .auto_in_awid(axi4index_auto_in_awid),
    .auto_in_awaddr(axi4index_auto_in_awaddr),
    .auto_in_awlen(axi4index_auto_in_awlen),
    .auto_in_awsize(axi4index_auto_in_awsize),
    .auto_in_awburst(axi4index_auto_in_awburst),
    .auto_in_awlock(axi4index_auto_in_awlock),
    .auto_in_awcache(axi4index_auto_in_awcache),
    .auto_in_awprot(axi4index_auto_in_awprot),
    .auto_in_awqos(axi4index_auto_in_awqos),
    .auto_in_awuser(axi4index_auto_in_awuser),
    .auto_in_awinstret(axi4index_auto_in_awinstret),
    .auto_in_wready(axi4index_auto_in_wready),
    .auto_in_wvalid(axi4index_auto_in_wvalid),
    .auto_in_wdata(axi4index_auto_in_wdata),
    .auto_in_wstrb(axi4index_auto_in_wstrb),
    .auto_in_wlast(axi4index_auto_in_wlast),
    .auto_in_bready(axi4index_auto_in_bready),
    .auto_in_bvalid(axi4index_auto_in_bvalid),
    .auto_in_bid(axi4index_auto_in_bid),
    .auto_in_bresp(axi4index_auto_in_bresp),
    .auto_in_buser(axi4index_auto_in_buser),
    .auto_in_arready(axi4index_auto_in_arready),
    .auto_in_arvalid(axi4index_auto_in_arvalid),
    .auto_in_arid(axi4index_auto_in_arid),
    .auto_in_araddr(axi4index_auto_in_araddr),
    .auto_in_arlen(axi4index_auto_in_arlen),
    .auto_in_arsize(axi4index_auto_in_arsize),
    .auto_in_arburst(axi4index_auto_in_arburst),
    .auto_in_arlock(axi4index_auto_in_arlock),
    .auto_in_arcache(axi4index_auto_in_arcache),
    .auto_in_arprot(axi4index_auto_in_arprot),
    .auto_in_arqos(axi4index_auto_in_arqos),
    .auto_in_aruser(axi4index_auto_in_aruser),
    .auto_in_arinstret(axi4index_auto_in_arinstret),
    .auto_in_rready(axi4index_auto_in_rready),
    .auto_in_rvalid(axi4index_auto_in_rvalid),
    .auto_in_rid(axi4index_auto_in_rid),
    .auto_in_rdata(axi4index_auto_in_rdata),
    .auto_in_rresp(axi4index_auto_in_rresp),
    .auto_in_ruser(axi4index_auto_in_ruser),
    .auto_in_rlast(axi4index_auto_in_rlast),
    .auto_out_awready(axi4index_auto_out_awready),
    .auto_out_awvalid(axi4index_auto_out_awvalid),
    .auto_out_awid(axi4index_auto_out_awid),
    .auto_out_awaddr(axi4index_auto_out_awaddr),
    .auto_out_awlen(axi4index_auto_out_awlen),
    .auto_out_awsize(axi4index_auto_out_awsize),
    .auto_out_awburst(axi4index_auto_out_awburst),
    .auto_out_awlock(axi4index_auto_out_awlock),
    .auto_out_awcache(axi4index_auto_out_awcache),
    .auto_out_awprot(axi4index_auto_out_awprot),
    .auto_out_awqos(axi4index_auto_out_awqos),
    .auto_out_awuser(axi4index_auto_out_awuser),
    .auto_out_awinstret(axi4index_auto_out_awinstret),
    .auto_out_wready(axi4index_auto_out_wready),
    .auto_out_wvalid(axi4index_auto_out_wvalid),
    .auto_out_wdata(axi4index_auto_out_wdata),
    .auto_out_wstrb(axi4index_auto_out_wstrb),
    .auto_out_wlast(axi4index_auto_out_wlast),
    .auto_out_bready(axi4index_auto_out_bready),
    .auto_out_bvalid(axi4index_auto_out_bvalid),
    .auto_out_bid(axi4index_auto_out_bid),
    .auto_out_bresp(axi4index_auto_out_bresp),
    .auto_out_buser(axi4index_auto_out_buser),
    .auto_out_arready(axi4index_auto_out_arready),
    .auto_out_arvalid(axi4index_auto_out_arvalid),
    .auto_out_arid(axi4index_auto_out_arid),
    .auto_out_araddr(axi4index_auto_out_araddr),
    .auto_out_arlen(axi4index_auto_out_arlen),
    .auto_out_arsize(axi4index_auto_out_arsize),
    .auto_out_arburst(axi4index_auto_out_arburst),
    .auto_out_arlock(axi4index_auto_out_arlock),
    .auto_out_arcache(axi4index_auto_out_arcache),
    .auto_out_arprot(axi4index_auto_out_arprot),
    .auto_out_arqos(axi4index_auto_out_arqos),
    .auto_out_aruser(axi4index_auto_out_aruser),
    .auto_out_arinstret(axi4index_auto_out_arinstret),
    .auto_out_rready(axi4index_auto_out_rready),
    .auto_out_rvalid(axi4index_auto_out_rvalid),
    .auto_out_rid(axi4index_auto_out_rid),
    .auto_out_rdata(axi4index_auto_out_rdata),
    .auto_out_rresp(axi4index_auto_out_rresp),
    .auto_out_ruser(axi4index_auto_out_ruser),
    .auto_out_rlast(axi4index_auto_out_rlast)
  );
  dual_TLToAXI4 tl2axi4 ( 
    .clock(tl2axi4_clock),
    .reset(tl2axi4_reset),
    .auto_in_a_ready(tl2axi4_auto_in_a_ready),
    .auto_in_a_valid(tl2axi4_auto_in_a_valid),
    .auto_in_a_bits_opcode(tl2axi4_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(tl2axi4_auto_in_a_bits_param),
    .auto_in_a_bits_size(tl2axi4_auto_in_a_bits_size),
    .auto_in_a_bits_source(tl2axi4_auto_in_a_bits_source),
    .auto_in_a_bits_address(tl2axi4_auto_in_a_bits_address),
    .auto_in_a_bits_mask(tl2axi4_auto_in_a_bits_mask),
    .auto_in_a_bits_data(tl2axi4_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(tl2axi4_auto_in_a_bits_corrupt),
    .auto_in_d_ready(tl2axi4_auto_in_d_ready),
    .auto_in_d_valid(tl2axi4_auto_in_d_valid),
    .auto_in_d_bits_opcode(tl2axi4_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(tl2axi4_auto_in_d_bits_size),
    .auto_in_d_bits_source(tl2axi4_auto_in_d_bits_source),
    .auto_in_d_bits_denied(tl2axi4_auto_in_d_bits_denied),
    .auto_in_d_bits_data(tl2axi4_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(tl2axi4_auto_in_d_bits_corrupt),
    .auto_out_awready(tl2axi4_auto_out_awready),
    .auto_out_awvalid(tl2axi4_auto_out_awvalid),
    .auto_out_awid(tl2axi4_auto_out_awid),
    .auto_out_awaddr(tl2axi4_auto_out_awaddr),
    .auto_out_awlen(tl2axi4_auto_out_awlen),
    .auto_out_awsize(tl2axi4_auto_out_awsize),
    .auto_out_awburst(tl2axi4_auto_out_awburst),
    .auto_out_awlock(tl2axi4_auto_out_awlock),
    .auto_out_awcache(tl2axi4_auto_out_awcache),
    .auto_out_awprot(tl2axi4_auto_out_awprot),
    .auto_out_awqos(tl2axi4_auto_out_awqos),
    .auto_out_awuser(tl2axi4_auto_out_awuser),
    .auto_out_awinstret(tl2axi4_auto_out_awinstret),
    .auto_out_wready(tl2axi4_auto_out_wready),
    .auto_out_wvalid(tl2axi4_auto_out_wvalid),
    .auto_out_wdata(tl2axi4_auto_out_wdata),
    .auto_out_wstrb(tl2axi4_auto_out_wstrb),
    .auto_out_wlast(tl2axi4_auto_out_wlast),
    .auto_out_bready(tl2axi4_auto_out_bready),
    .auto_out_bvalid(tl2axi4_auto_out_bvalid),
    .auto_out_bid(tl2axi4_auto_out_bid),
    .auto_out_bresp(tl2axi4_auto_out_bresp),
    .auto_out_buser(tl2axi4_auto_out_buser),
    .auto_out_arready(tl2axi4_auto_out_arready),
    .auto_out_arvalid(tl2axi4_auto_out_arvalid),
    .auto_out_arid(tl2axi4_auto_out_arid),
    .auto_out_araddr(tl2axi4_auto_out_araddr),
    .auto_out_arlen(tl2axi4_auto_out_arlen),
    .auto_out_arsize(tl2axi4_auto_out_arsize),
    .auto_out_arburst(tl2axi4_auto_out_arburst),
    .auto_out_arlock(tl2axi4_auto_out_arlock),
    .auto_out_arcache(tl2axi4_auto_out_arcache),
    .auto_out_arprot(tl2axi4_auto_out_arprot),
    .auto_out_arqos(tl2axi4_auto_out_arqos),
    .auto_out_aruser(tl2axi4_auto_out_aruser),
    .auto_out_arinstret(tl2axi4_auto_out_arinstret),
    .auto_out_rready(tl2axi4_auto_out_rready),
    .auto_out_rvalid(tl2axi4_auto_out_rvalid),
    .auto_out_rid(tl2axi4_auto_out_rid),
    .auto_out_rdata(tl2axi4_auto_out_rdata),
    .auto_out_rresp(tl2axi4_auto_out_rresp),
    .auto_out_ruser(tl2axi4_auto_out_ruser),
    .auto_out_rlast(tl2axi4_auto_out_rlast)
  );
  dual_AXI4Buffer axi4buf ( 
    .clock(axi4buf_clock),
    .reset(axi4buf_reset),
    .auto_in_awready(axi4buf_auto_in_awready),
    .auto_in_awvalid(axi4buf_auto_in_awvalid),
    .auto_in_awaddr(axi4buf_auto_in_awaddr),
    .auto_in_awlen(axi4buf_auto_in_awlen),
    .auto_in_awsize(axi4buf_auto_in_awsize),
    .auto_in_awburst(axi4buf_auto_in_awburst),
    .auto_in_awlock(axi4buf_auto_in_awlock),
    .auto_in_awcache(axi4buf_auto_in_awcache),
    .auto_in_awprot(axi4buf_auto_in_awprot),
    .auto_in_awqos(axi4buf_auto_in_awqos),
    .auto_in_awinstret(axi4buf_auto_in_awinstret),
    .auto_in_wready(axi4buf_auto_in_wready),
    .auto_in_wvalid(axi4buf_auto_in_wvalid),
    .auto_in_wdata(axi4buf_auto_in_wdata),
    .auto_in_wstrb(axi4buf_auto_in_wstrb),
    .auto_in_wlast(axi4buf_auto_in_wlast),
    .auto_in_bready(axi4buf_auto_in_bready),
    .auto_in_bvalid(axi4buf_auto_in_bvalid),
    .auto_in_bresp(axi4buf_auto_in_bresp),
    .auto_in_arready(axi4buf_auto_in_arready),
    .auto_in_arvalid(axi4buf_auto_in_arvalid),
    .auto_in_araddr(axi4buf_auto_in_araddr),
    .auto_in_arlen(axi4buf_auto_in_arlen),
    .auto_in_arsize(axi4buf_auto_in_arsize),
    .auto_in_arburst(axi4buf_auto_in_arburst),
    .auto_in_arlock(axi4buf_auto_in_arlock),
    .auto_in_arcache(axi4buf_auto_in_arcache),
    .auto_in_arprot(axi4buf_auto_in_arprot),
    .auto_in_arqos(axi4buf_auto_in_arqos),
    .auto_in_arinstret(axi4buf_auto_in_arinstret),
    .auto_in_rready(axi4buf_auto_in_rready),
    .auto_in_rvalid(axi4buf_auto_in_rvalid),
    .auto_in_rdata(axi4buf_auto_in_rdata),
    .auto_in_rresp(axi4buf_auto_in_rresp),
    .auto_in_rlast(axi4buf_auto_in_rlast),
    .auto_out_awready(axi4buf_auto_out_awready),
    .auto_out_awvalid(axi4buf_auto_out_awvalid),
    .auto_out_awid(axi4buf_auto_out_awid),
    .auto_out_awaddr(axi4buf_auto_out_awaddr),
    .auto_out_awlen(axi4buf_auto_out_awlen),
    .auto_out_awsize(axi4buf_auto_out_awsize),
    .auto_out_awburst(axi4buf_auto_out_awburst),
    .auto_out_awlock(axi4buf_auto_out_awlock),
    .auto_out_awcache(axi4buf_auto_out_awcache),
    .auto_out_awprot(axi4buf_auto_out_awprot),
    .auto_out_awqos(axi4buf_auto_out_awqos),
    .auto_out_awinstret(axi4buf_auto_out_awinstret),
    .auto_out_wready(axi4buf_auto_out_wready),
    .auto_out_wvalid(axi4buf_auto_out_wvalid),
    .auto_out_wdata(axi4buf_auto_out_wdata),
    .auto_out_wstrb(axi4buf_auto_out_wstrb),
    .auto_out_wlast(axi4buf_auto_out_wlast),
    .auto_out_bready(axi4buf_auto_out_bready),
    .auto_out_bvalid(axi4buf_auto_out_bvalid),
    .auto_out_bresp(axi4buf_auto_out_bresp),
    .auto_out_arready(axi4buf_auto_out_arready),
    .auto_out_arvalid(axi4buf_auto_out_arvalid),
    .auto_out_arid(axi4buf_auto_out_arid),
    .auto_out_araddr(axi4buf_auto_out_araddr),
    .auto_out_arlen(axi4buf_auto_out_arlen),
    .auto_out_arsize(axi4buf_auto_out_arsize),
    .auto_out_arburst(axi4buf_auto_out_arburst),
    .auto_out_arlock(axi4buf_auto_out_arlock),
    .auto_out_arcache(axi4buf_auto_out_arcache),
    .auto_out_arprot(axi4buf_auto_out_arprot),
    .auto_out_arqos(axi4buf_auto_out_arqos),
    .auto_out_arinstret(axi4buf_auto_out_arinstret),
    .auto_out_rready(axi4buf_auto_out_rready),
    .auto_out_rvalid(axi4buf_auto_out_rvalid),
    .auto_out_rdata(axi4buf_auto_out_rdata),
    .auto_out_rresp(axi4buf_auto_out_rresp),
    .auto_out_rlast(axi4buf_auto_out_rlast)
  );
  dual_AXI4UserYanker_1 axi4yank_1 ( 
    .clock(axi4yank_1_clock),
    .reset(axi4yank_1_reset),
    .auto_in_awready(axi4yank_1_auto_in_awready),
    .auto_in_awvalid(axi4yank_1_auto_in_awvalid),
    .auto_in_awaddr(axi4yank_1_auto_in_awaddr),
    .auto_in_awlen(axi4yank_1_auto_in_awlen),
    .auto_in_awsize(axi4yank_1_auto_in_awsize),
    .auto_in_awburst(axi4yank_1_auto_in_awburst),
    .auto_in_awlock(axi4yank_1_auto_in_awlock),
    .auto_in_awcache(axi4yank_1_auto_in_awcache),
    .auto_in_awprot(axi4yank_1_auto_in_awprot),
    .auto_in_awqos(axi4yank_1_auto_in_awqos),
    .auto_in_awuser(axi4yank_1_auto_in_awuser),
    .auto_in_awinstret(axi4yank_1_auto_in_awinstret),
    .auto_in_wready(axi4yank_1_auto_in_wready),
    .auto_in_wvalid(axi4yank_1_auto_in_wvalid),
    .auto_in_wdata(axi4yank_1_auto_in_wdata),
    .auto_in_wstrb(axi4yank_1_auto_in_wstrb),
    .auto_in_wlast(axi4yank_1_auto_in_wlast),
    .auto_in_bready(axi4yank_1_auto_in_bready),
    .auto_in_bvalid(axi4yank_1_auto_in_bvalid),
    .auto_in_bresp(axi4yank_1_auto_in_bresp),
    .auto_in_buser(axi4yank_1_auto_in_buser),
    .auto_in_arready(axi4yank_1_auto_in_arready),
    .auto_in_arvalid(axi4yank_1_auto_in_arvalid),
    .auto_in_araddr(axi4yank_1_auto_in_araddr),
    .auto_in_arlen(axi4yank_1_auto_in_arlen),
    .auto_in_arsize(axi4yank_1_auto_in_arsize),
    .auto_in_arburst(axi4yank_1_auto_in_arburst),
    .auto_in_arlock(axi4yank_1_auto_in_arlock),
    .auto_in_arcache(axi4yank_1_auto_in_arcache),
    .auto_in_arprot(axi4yank_1_auto_in_arprot),
    .auto_in_arqos(axi4yank_1_auto_in_arqos),
    .auto_in_aruser(axi4yank_1_auto_in_aruser),
    .auto_in_arinstret(axi4yank_1_auto_in_arinstret),
    .auto_in_rready(axi4yank_1_auto_in_rready),
    .auto_in_rvalid(axi4yank_1_auto_in_rvalid),
    .auto_in_rdata(axi4yank_1_auto_in_rdata),
    .auto_in_rresp(axi4yank_1_auto_in_rresp),
    .auto_in_ruser(axi4yank_1_auto_in_ruser),
    .auto_in_rlast(axi4yank_1_auto_in_rlast),
    .auto_out_awready(axi4yank_1_auto_out_awready),
    .auto_out_awvalid(axi4yank_1_auto_out_awvalid),
    .auto_out_awaddr(axi4yank_1_auto_out_awaddr),
    .auto_out_awlen(axi4yank_1_auto_out_awlen),
    .auto_out_awsize(axi4yank_1_auto_out_awsize),
    .auto_out_awburst(axi4yank_1_auto_out_awburst),
    .auto_out_awlock(axi4yank_1_auto_out_awlock),
    .auto_out_awcache(axi4yank_1_auto_out_awcache),
    .auto_out_awprot(axi4yank_1_auto_out_awprot),
    .auto_out_awqos(axi4yank_1_auto_out_awqos),
    .auto_out_awinstret(axi4yank_1_auto_out_awinstret),
    .auto_out_wready(axi4yank_1_auto_out_wready),
    .auto_out_wvalid(axi4yank_1_auto_out_wvalid),
    .auto_out_wdata(axi4yank_1_auto_out_wdata),
    .auto_out_wstrb(axi4yank_1_auto_out_wstrb),
    .auto_out_wlast(axi4yank_1_auto_out_wlast),
    .auto_out_bready(axi4yank_1_auto_out_bready),
    .auto_out_bvalid(axi4yank_1_auto_out_bvalid),
    .auto_out_bresp(axi4yank_1_auto_out_bresp),
    .auto_out_arready(axi4yank_1_auto_out_arready),
    .auto_out_arvalid(axi4yank_1_auto_out_arvalid),
    .auto_out_araddr(axi4yank_1_auto_out_araddr),
    .auto_out_arlen(axi4yank_1_auto_out_arlen),
    .auto_out_arsize(axi4yank_1_auto_out_arsize),
    .auto_out_arburst(axi4yank_1_auto_out_arburst),
    .auto_out_arlock(axi4yank_1_auto_out_arlock),
    .auto_out_arcache(axi4yank_1_auto_out_arcache),
    .auto_out_arprot(axi4yank_1_auto_out_arprot),
    .auto_out_arqos(axi4yank_1_auto_out_arqos),
    .auto_out_arinstret(axi4yank_1_auto_out_arinstret),
    .auto_out_rready(axi4yank_1_auto_out_rready),
    .auto_out_rvalid(axi4yank_1_auto_out_rvalid),
    .auto_out_rdata(axi4yank_1_auto_out_rdata),
    .auto_out_rresp(axi4yank_1_auto_out_rresp),
    .auto_out_rlast(axi4yank_1_auto_out_rlast)
  );
  dual_AXI4Deinterleaver axi4deint ( 
    .clock(axi4deint_clock),
    .reset(axi4deint_reset),
    .auto_in_awready(axi4deint_auto_in_awready),
    .auto_in_awvalid(axi4deint_auto_in_awvalid),
    .auto_in_awaddr(axi4deint_auto_in_awaddr),
    .auto_in_awlen(axi4deint_auto_in_awlen),
    .auto_in_awsize(axi4deint_auto_in_awsize),
    .auto_in_awburst(axi4deint_auto_in_awburst),
    .auto_in_awlock(axi4deint_auto_in_awlock),
    .auto_in_awcache(axi4deint_auto_in_awcache),
    .auto_in_awprot(axi4deint_auto_in_awprot),
    .auto_in_awqos(axi4deint_auto_in_awqos),
    .auto_in_awuser(axi4deint_auto_in_awuser),
    .auto_in_awinstret(axi4deint_auto_in_awinstret),
    .auto_in_wready(axi4deint_auto_in_wready),
    .auto_in_wvalid(axi4deint_auto_in_wvalid),
    .auto_in_wdata(axi4deint_auto_in_wdata),
    .auto_in_wstrb(axi4deint_auto_in_wstrb),
    .auto_in_wlast(axi4deint_auto_in_wlast),
    .auto_in_bready(axi4deint_auto_in_bready),
    .auto_in_bvalid(axi4deint_auto_in_bvalid),
    .auto_in_bresp(axi4deint_auto_in_bresp),
    .auto_in_buser(axi4deint_auto_in_buser),
    .auto_in_arready(axi4deint_auto_in_arready),
    .auto_in_arvalid(axi4deint_auto_in_arvalid),
    .auto_in_araddr(axi4deint_auto_in_araddr),
    .auto_in_arlen(axi4deint_auto_in_arlen),
    .auto_in_arsize(axi4deint_auto_in_arsize),
    .auto_in_arburst(axi4deint_auto_in_arburst),
    .auto_in_arlock(axi4deint_auto_in_arlock),
    .auto_in_arcache(axi4deint_auto_in_arcache),
    .auto_in_arprot(axi4deint_auto_in_arprot),
    .auto_in_arqos(axi4deint_auto_in_arqos),
    .auto_in_aruser(axi4deint_auto_in_aruser),
    .auto_in_arinstret(axi4deint_auto_in_arinstret),
    .auto_in_rready(axi4deint_auto_in_rready),
    .auto_in_rvalid(axi4deint_auto_in_rvalid),
    .auto_in_rdata(axi4deint_auto_in_rdata),
    .auto_in_rresp(axi4deint_auto_in_rresp),
    .auto_in_ruser(axi4deint_auto_in_ruser),
    .auto_in_rlast(axi4deint_auto_in_rlast),
    .auto_out_awready(axi4deint_auto_out_awready),
    .auto_out_awvalid(axi4deint_auto_out_awvalid),
    .auto_out_awaddr(axi4deint_auto_out_awaddr),
    .auto_out_awlen(axi4deint_auto_out_awlen),
    .auto_out_awsize(axi4deint_auto_out_awsize),
    .auto_out_awburst(axi4deint_auto_out_awburst),
    .auto_out_awlock(axi4deint_auto_out_awlock),
    .auto_out_awcache(axi4deint_auto_out_awcache),
    .auto_out_awprot(axi4deint_auto_out_awprot),
    .auto_out_awqos(axi4deint_auto_out_awqos),
    .auto_out_awuser(axi4deint_auto_out_awuser),
    .auto_out_awinstret(axi4deint_auto_out_awinstret),
    .auto_out_wready(axi4deint_auto_out_wready),
    .auto_out_wvalid(axi4deint_auto_out_wvalid),
    .auto_out_wdata(axi4deint_auto_out_wdata),
    .auto_out_wstrb(axi4deint_auto_out_wstrb),
    .auto_out_wlast(axi4deint_auto_out_wlast),
    .auto_out_bready(axi4deint_auto_out_bready),
    .auto_out_bvalid(axi4deint_auto_out_bvalid),
    .auto_out_bresp(axi4deint_auto_out_bresp),
    .auto_out_buser(axi4deint_auto_out_buser),
    .auto_out_arready(axi4deint_auto_out_arready),
    .auto_out_arvalid(axi4deint_auto_out_arvalid),
    .auto_out_araddr(axi4deint_auto_out_araddr),
    .auto_out_arlen(axi4deint_auto_out_arlen),
    .auto_out_arsize(axi4deint_auto_out_arsize),
    .auto_out_arburst(axi4deint_auto_out_arburst),
    .auto_out_arlock(axi4deint_auto_out_arlock),
    .auto_out_arcache(axi4deint_auto_out_arcache),
    .auto_out_arprot(axi4deint_auto_out_arprot),
    .auto_out_arqos(axi4deint_auto_out_arqos),
    .auto_out_aruser(axi4deint_auto_out_aruser),
    .auto_out_arinstret(axi4deint_auto_out_arinstret),
    .auto_out_rready(axi4deint_auto_out_rready),
    .auto_out_rvalid(axi4deint_auto_out_rvalid),
    .auto_out_rdata(axi4deint_auto_out_rdata),
    .auto_out_rresp(axi4deint_auto_out_rresp),
    .auto_out_ruser(axi4deint_auto_out_ruser),
    .auto_out_rlast(axi4deint_auto_out_rlast)
  );
  dual_AXI4IdIndexer_1 axi4index_1 ( 
    .auto_in_awready(axi4index_1_auto_in_awready),
    .auto_in_awvalid(axi4index_1_auto_in_awvalid),
    .auto_in_awid(axi4index_1_auto_in_awid),
    .auto_in_awaddr(axi4index_1_auto_in_awaddr),
    .auto_in_awlen(axi4index_1_auto_in_awlen),
    .auto_in_awsize(axi4index_1_auto_in_awsize),
    .auto_in_awburst(axi4index_1_auto_in_awburst),
    .auto_in_awlock(axi4index_1_auto_in_awlock),
    .auto_in_awcache(axi4index_1_auto_in_awcache),
    .auto_in_awprot(axi4index_1_auto_in_awprot),
    .auto_in_awqos(axi4index_1_auto_in_awqos),
    .auto_in_awuser(axi4index_1_auto_in_awuser),
    .auto_in_awinstret(axi4index_1_auto_in_awinstret),
    .auto_in_wready(axi4index_1_auto_in_wready),
    .auto_in_wvalid(axi4index_1_auto_in_wvalid),
    .auto_in_wdata(axi4index_1_auto_in_wdata),
    .auto_in_wstrb(axi4index_1_auto_in_wstrb),
    .auto_in_wlast(axi4index_1_auto_in_wlast),
    .auto_in_bready(axi4index_1_auto_in_bready),
    .auto_in_bvalid(axi4index_1_auto_in_bvalid),
    .auto_in_bid(axi4index_1_auto_in_bid),
    .auto_in_bresp(axi4index_1_auto_in_bresp),
    .auto_in_buser(axi4index_1_auto_in_buser),
    .auto_in_arready(axi4index_1_auto_in_arready),
    .auto_in_arvalid(axi4index_1_auto_in_arvalid),
    .auto_in_arid(axi4index_1_auto_in_arid),
    .auto_in_araddr(axi4index_1_auto_in_araddr),
    .auto_in_arlen(axi4index_1_auto_in_arlen),
    .auto_in_arsize(axi4index_1_auto_in_arsize),
    .auto_in_arburst(axi4index_1_auto_in_arburst),
    .auto_in_arlock(axi4index_1_auto_in_arlock),
    .auto_in_arcache(axi4index_1_auto_in_arcache),
    .auto_in_arprot(axi4index_1_auto_in_arprot),
    .auto_in_arqos(axi4index_1_auto_in_arqos),
    .auto_in_aruser(axi4index_1_auto_in_aruser),
    .auto_in_arinstret(axi4index_1_auto_in_arinstret),
    .auto_in_rready(axi4index_1_auto_in_rready),
    .auto_in_rvalid(axi4index_1_auto_in_rvalid),
    .auto_in_rid(axi4index_1_auto_in_rid),
    .auto_in_rdata(axi4index_1_auto_in_rdata),
    .auto_in_rresp(axi4index_1_auto_in_rresp),
    .auto_in_ruser(axi4index_1_auto_in_ruser),
    .auto_in_rlast(axi4index_1_auto_in_rlast),
    .auto_out_awready(axi4index_1_auto_out_awready),
    .auto_out_awvalid(axi4index_1_auto_out_awvalid),
    .auto_out_awaddr(axi4index_1_auto_out_awaddr),
    .auto_out_awlen(axi4index_1_auto_out_awlen),
    .auto_out_awsize(axi4index_1_auto_out_awsize),
    .auto_out_awburst(axi4index_1_auto_out_awburst),
    .auto_out_awlock(axi4index_1_auto_out_awlock),
    .auto_out_awcache(axi4index_1_auto_out_awcache),
    .auto_out_awprot(axi4index_1_auto_out_awprot),
    .auto_out_awqos(axi4index_1_auto_out_awqos),
    .auto_out_awuser(axi4index_1_auto_out_awuser),
    .auto_out_awinstret(axi4index_1_auto_out_awinstret),
    .auto_out_wready(axi4index_1_auto_out_wready),
    .auto_out_wvalid(axi4index_1_auto_out_wvalid),
    .auto_out_wdata(axi4index_1_auto_out_wdata),
    .auto_out_wstrb(axi4index_1_auto_out_wstrb),
    .auto_out_wlast(axi4index_1_auto_out_wlast),
    .auto_out_bready(axi4index_1_auto_out_bready),
    .auto_out_bvalid(axi4index_1_auto_out_bvalid),
    .auto_out_bresp(axi4index_1_auto_out_bresp),
    .auto_out_buser(axi4index_1_auto_out_buser),
    .auto_out_arready(axi4index_1_auto_out_arready),
    .auto_out_arvalid(axi4index_1_auto_out_arvalid),
    .auto_out_araddr(axi4index_1_auto_out_araddr),
    .auto_out_arlen(axi4index_1_auto_out_arlen),
    .auto_out_arsize(axi4index_1_auto_out_arsize),
    .auto_out_arburst(axi4index_1_auto_out_arburst),
    .auto_out_arlock(axi4index_1_auto_out_arlock),
    .auto_out_arcache(axi4index_1_auto_out_arcache),
    .auto_out_arprot(axi4index_1_auto_out_arprot),
    .auto_out_arqos(axi4index_1_auto_out_arqos),
    .auto_out_aruser(axi4index_1_auto_out_aruser),
    .auto_out_arinstret(axi4index_1_auto_out_arinstret),
    .auto_out_rready(axi4index_1_auto_out_rready),
    .auto_out_rvalid(axi4index_1_auto_out_rvalid),
    .auto_out_rdata(axi4index_1_auto_out_rdata),
    .auto_out_rresp(axi4index_1_auto_out_rresp),
    .auto_out_ruser(axi4index_1_auto_out_ruser),
    .auto_out_rlast(axi4index_1_auto_out_rlast)
  );
  dual_TLToAXI4_1 tl2axi4_1 ( 
    .clock(tl2axi4_1_clock),
    .reset(tl2axi4_1_reset),
    .auto_in_a_ready(tl2axi4_1_auto_in_a_ready),
    .auto_in_a_valid(tl2axi4_1_auto_in_a_valid),
    .auto_in_a_bits_opcode(tl2axi4_1_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(tl2axi4_1_auto_in_a_bits_param),
    .auto_in_a_bits_size(tl2axi4_1_auto_in_a_bits_size),
    .auto_in_a_bits_source(tl2axi4_1_auto_in_a_bits_source),
    .auto_in_a_bits_address(tl2axi4_1_auto_in_a_bits_address),
    .auto_in_a_bits_mask(tl2axi4_1_auto_in_a_bits_mask),
    .auto_in_a_bits_data(tl2axi4_1_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(tl2axi4_1_auto_in_a_bits_corrupt),
    .auto_in_d_ready(tl2axi4_1_auto_in_d_ready),
    .auto_in_d_valid(tl2axi4_1_auto_in_d_valid),
    .auto_in_d_bits_opcode(tl2axi4_1_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(tl2axi4_1_auto_in_d_bits_size),
    .auto_in_d_bits_source(tl2axi4_1_auto_in_d_bits_source),
    .auto_in_d_bits_denied(tl2axi4_1_auto_in_d_bits_denied),
    .auto_in_d_bits_data(tl2axi4_1_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(tl2axi4_1_auto_in_d_bits_corrupt),
    .auto_out_awready(tl2axi4_1_auto_out_awready),
    .auto_out_awvalid(tl2axi4_1_auto_out_awvalid),
    .auto_out_awid(tl2axi4_1_auto_out_awid),
    .auto_out_awaddr(tl2axi4_1_auto_out_awaddr),
    .auto_out_awlen(tl2axi4_1_auto_out_awlen),
    .auto_out_awsize(tl2axi4_1_auto_out_awsize),
    .auto_out_awburst(tl2axi4_1_auto_out_awburst),
    .auto_out_awlock(tl2axi4_1_auto_out_awlock),
    .auto_out_awcache(tl2axi4_1_auto_out_awcache),
    .auto_out_awprot(tl2axi4_1_auto_out_awprot),
    .auto_out_awqos(tl2axi4_1_auto_out_awqos),
    .auto_out_awuser(tl2axi4_1_auto_out_awuser),
    .auto_out_awinstret(tl2axi4_1_auto_out_awinstret),
    .auto_out_wready(tl2axi4_1_auto_out_wready),
    .auto_out_wvalid(tl2axi4_1_auto_out_wvalid),
    .auto_out_wdata(tl2axi4_1_auto_out_wdata),
    .auto_out_wstrb(tl2axi4_1_auto_out_wstrb),
    .auto_out_wlast(tl2axi4_1_auto_out_wlast),
    .auto_out_bready(tl2axi4_1_auto_out_bready),
    .auto_out_bvalid(tl2axi4_1_auto_out_bvalid),
    .auto_out_bid(tl2axi4_1_auto_out_bid),
    .auto_out_bresp(tl2axi4_1_auto_out_bresp),
    .auto_out_buser(tl2axi4_1_auto_out_buser),
    .auto_out_arready(tl2axi4_1_auto_out_arready),
    .auto_out_arvalid(tl2axi4_1_auto_out_arvalid),
    .auto_out_arid(tl2axi4_1_auto_out_arid),
    .auto_out_araddr(tl2axi4_1_auto_out_araddr),
    .auto_out_arlen(tl2axi4_1_auto_out_arlen),
    .auto_out_arsize(tl2axi4_1_auto_out_arsize),
    .auto_out_arburst(tl2axi4_1_auto_out_arburst),
    .auto_out_arlock(tl2axi4_1_auto_out_arlock),
    .auto_out_arcache(tl2axi4_1_auto_out_arcache),
    .auto_out_arprot(tl2axi4_1_auto_out_arprot),
    .auto_out_arqos(tl2axi4_1_auto_out_arqos),
    .auto_out_aruser(tl2axi4_1_auto_out_aruser),
    .auto_out_arinstret(tl2axi4_1_auto_out_arinstret),
    .auto_out_rready(tl2axi4_1_auto_out_rready),
    .auto_out_rvalid(tl2axi4_1_auto_out_rvalid),
    .auto_out_rid(tl2axi4_1_auto_out_rid),
    .auto_out_rdata(tl2axi4_1_auto_out_rdata),
    .auto_out_rresp(tl2axi4_1_auto_out_rresp),
    .auto_out_ruser(tl2axi4_1_auto_out_ruser),
    .auto_out_rlast(tl2axi4_1_auto_out_rlast)
  );
  dual_TLFIFOFixer fixer ( 
    .clock(fixer_clock),
    .reset(fixer_reset),
    .auto_in_a_ready(fixer_auto_in_a_ready),
    .auto_in_a_valid(fixer_auto_in_a_valid),
    .auto_in_a_bits_opcode(fixer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(fixer_auto_in_a_bits_param),
    .auto_in_a_bits_size(fixer_auto_in_a_bits_size),
    .auto_in_a_bits_source(fixer_auto_in_a_bits_source),
    .auto_in_a_bits_address(fixer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fixer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(fixer_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(fixer_auto_in_a_bits_corrupt),
    .auto_in_d_ready(fixer_auto_in_d_ready),
    .auto_in_d_valid(fixer_auto_in_d_valid),
    .auto_in_d_bits_opcode(fixer_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(fixer_auto_in_d_bits_param),
    .auto_in_d_bits_size(fixer_auto_in_d_bits_size),
    .auto_in_d_bits_source(fixer_auto_in_d_bits_source),
    .auto_in_d_bits_sink(fixer_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(fixer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(fixer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(fixer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(fixer_auto_out_a_ready),
    .auto_out_a_valid(fixer_auto_out_a_valid),
    .auto_out_a_bits_opcode(fixer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(fixer_auto_out_a_bits_param),
    .auto_out_a_bits_size(fixer_auto_out_a_bits_size),
    .auto_out_a_bits_source(fixer_auto_out_a_bits_source),
    .auto_out_a_bits_address(fixer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(fixer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(fixer_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(fixer_auto_out_a_bits_corrupt),
    .auto_out_d_ready(fixer_auto_out_d_ready),
    .auto_out_d_valid(fixer_auto_out_d_valid),
    .auto_out_d_bits_opcode(fixer_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(fixer_auto_out_d_bits_param),
    .auto_out_d_bits_size(fixer_auto_out_d_bits_size),
    .auto_out_d_bits_source(fixer_auto_out_d_bits_source),
    .auto_out_d_bits_sink(fixer_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(fixer_auto_out_d_bits_denied),
    .auto_out_d_bits_data(fixer_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(fixer_auto_out_d_bits_corrupt)
  );
  dual_TLWidthWidget widget ( 
    .clock(widget_clock),
    .reset(widget_reset),
    .auto_in_a_ready(widget_auto_in_a_ready),
    .auto_in_a_valid(widget_auto_in_a_valid),
    .auto_in_a_bits_opcode(widget_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(widget_auto_in_a_bits_param),
    .auto_in_a_bits_size(widget_auto_in_a_bits_size),
    .auto_in_a_bits_source(widget_auto_in_a_bits_source),
    .auto_in_a_bits_address(widget_auto_in_a_bits_address),
    .auto_in_a_bits_mask(widget_auto_in_a_bits_mask),
    .auto_in_a_bits_data(widget_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(widget_auto_in_a_bits_corrupt),
    .auto_in_d_ready(widget_auto_in_d_ready),
    .auto_in_d_valid(widget_auto_in_d_valid),
    .auto_in_d_bits_opcode(widget_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(widget_auto_in_d_bits_size),
    .auto_in_d_bits_source(widget_auto_in_d_bits_source),
    .auto_in_d_bits_denied(widget_auto_in_d_bits_denied),
    .auto_in_d_bits_data(widget_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(widget_auto_in_d_bits_corrupt),
    .auto_out_a_ready(widget_auto_out_a_ready),
    .auto_out_a_valid(widget_auto_out_a_valid),
    .auto_out_a_bits_opcode(widget_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(widget_auto_out_a_bits_param),
    .auto_out_a_bits_size(widget_auto_out_a_bits_size),
    .auto_out_a_bits_source(widget_auto_out_a_bits_source),
    .auto_out_a_bits_address(widget_auto_out_a_bits_address),
    .auto_out_a_bits_mask(widget_auto_out_a_bits_mask),
    .auto_out_a_bits_data(widget_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(widget_auto_out_a_bits_corrupt),
    .auto_out_d_ready(widget_auto_out_d_ready),
    .auto_out_d_valid(widget_auto_out_d_valid),
    .auto_out_d_bits_opcode(widget_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(widget_auto_out_d_bits_param),
    .auto_out_d_bits_size(widget_auto_out_d_bits_size),
    .auto_out_d_bits_source(widget_auto_out_d_bits_source),
    .auto_out_d_bits_sink(widget_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(widget_auto_out_d_bits_denied),
    .auto_out_d_bits_data(widget_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(widget_auto_out_d_bits_corrupt)
  );
  dual_AXI4ToTL_top axi42tl ( 
    .clock(axi42tl_clock),
    .reset(axi42tl_reset),
    .auto_in_awready(axi42tl_auto_in_awready),
    .auto_in_awvalid(axi42tl_auto_in_awvalid),
    .auto_in_awid(axi42tl_auto_in_awid),
    .auto_in_awaddr(axi42tl_auto_in_awaddr),
    .auto_in_awlen(axi42tl_auto_in_awlen),
    .auto_in_awsize(axi42tl_auto_in_awsize),
    .auto_in_wready(axi42tl_auto_in_wready),
    .auto_in_wvalid(axi42tl_auto_in_wvalid),
    .auto_in_wdata(axi42tl_auto_in_wdata),
    .auto_in_wstrb(axi42tl_auto_in_wstrb),
    .auto_in_wlast(axi42tl_auto_in_wlast),
    .auto_in_bready(axi42tl_auto_in_bready),
    .auto_in_bvalid(axi42tl_auto_in_bvalid),
    .auto_in_bid(axi42tl_auto_in_bid),
    .auto_in_bresp(axi42tl_auto_in_bresp),
    .auto_in_arready(axi42tl_auto_in_arready),
    .auto_in_arvalid(axi42tl_auto_in_arvalid),
    .auto_in_arid(axi42tl_auto_in_arid),
    .auto_in_araddr(axi42tl_auto_in_araddr),
    .auto_in_arlen(axi42tl_auto_in_arlen),
    .auto_in_arsize(axi42tl_auto_in_arsize),
    .auto_in_rready(axi42tl_auto_in_rready),
    .auto_in_rvalid(axi42tl_auto_in_rvalid),
    .auto_in_rid(axi42tl_auto_in_rid),
    .auto_in_rdata(axi42tl_auto_in_rdata),
    .auto_in_rresp(axi42tl_auto_in_rresp),
    .auto_in_rlast(axi42tl_auto_in_rlast),
    .auto_out_a_ready(axi42tl_auto_out_a_ready),
    .auto_out_a_valid(axi42tl_auto_out_a_valid),
    .auto_out_a_bits_opcode(axi42tl_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(axi42tl_auto_out_a_bits_param),
    .auto_out_a_bits_size(axi42tl_auto_out_a_bits_size),
    .auto_out_a_bits_source(axi42tl_auto_out_a_bits_source),
    .auto_out_a_bits_address(axi42tl_auto_out_a_bits_address),
    .auto_out_a_bits_mask(axi42tl_auto_out_a_bits_mask),
    .auto_out_a_bits_data(axi42tl_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(axi42tl_auto_out_a_bits_corrupt),
    .auto_out_d_ready(axi42tl_auto_out_d_ready),
    .auto_out_d_valid(axi42tl_auto_out_d_valid),
    .auto_out_d_bits_opcode(axi42tl_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(axi42tl_auto_out_d_bits_size),
    .auto_out_d_bits_source(axi42tl_auto_out_d_bits_source),
    .auto_out_d_bits_denied(axi42tl_auto_out_d_bits_denied),
    .auto_out_d_bits_data(axi42tl_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(axi42tl_auto_out_d_bits_corrupt)
  );
  dual_AXI4UserYanker_2 axi4yank_2 ( 
    .clock(axi4yank_2_clock),
    .reset(axi4yank_2_reset),
    .auto_in_awready(axi4yank_2_auto_in_awready),
    .auto_in_awvalid(axi4yank_2_auto_in_awvalid),
    .auto_in_awid(axi4yank_2_auto_in_awid),
    .auto_in_awaddr(axi4yank_2_auto_in_awaddr),
    .auto_in_awlen(axi4yank_2_auto_in_awlen),
    .auto_in_awsize(axi4yank_2_auto_in_awsize),
    .auto_in_awuser(axi4yank_2_auto_in_awuser),
    .auto_in_wready(axi4yank_2_auto_in_wready),
    .auto_in_wvalid(axi4yank_2_auto_in_wvalid),
    .auto_in_wdata(axi4yank_2_auto_in_wdata),
    .auto_in_wstrb(axi4yank_2_auto_in_wstrb),
    .auto_in_wlast(axi4yank_2_auto_in_wlast),
    .auto_in_bready(axi4yank_2_auto_in_bready),
    .auto_in_bvalid(axi4yank_2_auto_in_bvalid),
    .auto_in_bid(axi4yank_2_auto_in_bid),
    .auto_in_bresp(axi4yank_2_auto_in_bresp),
    .auto_in_buser(axi4yank_2_auto_in_buser),
    .auto_in_arready(axi4yank_2_auto_in_arready),
    .auto_in_arvalid(axi4yank_2_auto_in_arvalid),
    .auto_in_arid(axi4yank_2_auto_in_arid),
    .auto_in_araddr(axi4yank_2_auto_in_araddr),
    .auto_in_arlen(axi4yank_2_auto_in_arlen),
    .auto_in_arsize(axi4yank_2_auto_in_arsize),
    .auto_in_aruser(axi4yank_2_auto_in_aruser),
    .auto_in_rready(axi4yank_2_auto_in_rready),
    .auto_in_rvalid(axi4yank_2_auto_in_rvalid),
    .auto_in_rid(axi4yank_2_auto_in_rid),
    .auto_in_rdata(axi4yank_2_auto_in_rdata),
    .auto_in_rresp(axi4yank_2_auto_in_rresp),
    .auto_in_ruser(axi4yank_2_auto_in_ruser),
    .auto_in_rlast(axi4yank_2_auto_in_rlast),
    .auto_out_awready(axi4yank_2_auto_out_awready),
    .auto_out_awvalid(axi4yank_2_auto_out_awvalid),
    .auto_out_awid(axi4yank_2_auto_out_awid),
    .auto_out_awaddr(axi4yank_2_auto_out_awaddr),
    .auto_out_awlen(axi4yank_2_auto_out_awlen),
    .auto_out_awsize(axi4yank_2_auto_out_awsize),
    .auto_out_wready(axi4yank_2_auto_out_wready),
    .auto_out_wvalid(axi4yank_2_auto_out_wvalid),
    .auto_out_wdata(axi4yank_2_auto_out_wdata),
    .auto_out_wstrb(axi4yank_2_auto_out_wstrb),
    .auto_out_wlast(axi4yank_2_auto_out_wlast),
    .auto_out_bready(axi4yank_2_auto_out_bready),
    .auto_out_bvalid(axi4yank_2_auto_out_bvalid),
    .auto_out_bid(axi4yank_2_auto_out_bid),
    .auto_out_bresp(axi4yank_2_auto_out_bresp),
    .auto_out_arready(axi4yank_2_auto_out_arready),
    .auto_out_arvalid(axi4yank_2_auto_out_arvalid),
    .auto_out_arid(axi4yank_2_auto_out_arid),
    .auto_out_araddr(axi4yank_2_auto_out_araddr),
    .auto_out_arlen(axi4yank_2_auto_out_arlen),
    .auto_out_arsize(axi4yank_2_auto_out_arsize),
    .auto_out_rready(axi4yank_2_auto_out_rready),
    .auto_out_rvalid(axi4yank_2_auto_out_rvalid),
    .auto_out_rid(axi4yank_2_auto_out_rid),
    .auto_out_rdata(axi4yank_2_auto_out_rdata),
    .auto_out_rresp(axi4yank_2_auto_out_rresp),
    .auto_out_rlast(axi4yank_2_auto_out_rlast)
  );
  dual_AXI4Fragmenter axi4frag ( 
    .clock(axi4frag_clock),
    .reset(axi4frag_reset),
    .auto_in_awready(axi4frag_auto_in_awready),
    .auto_in_awvalid(axi4frag_auto_in_awvalid),
    .auto_in_awid(axi4frag_auto_in_awid),
    .auto_in_awaddr(axi4frag_auto_in_awaddr),
    .auto_in_awlen(axi4frag_auto_in_awlen),
    .auto_in_awsize(axi4frag_auto_in_awsize),
    .auto_in_awburst(axi4frag_auto_in_awburst),
    .auto_in_awuser(axi4frag_auto_in_awuser),
    .auto_in_wready(axi4frag_auto_in_wready),
    .auto_in_wvalid(axi4frag_auto_in_wvalid),
    .auto_in_wdata(axi4frag_auto_in_wdata),
    .auto_in_wstrb(axi4frag_auto_in_wstrb),
    .auto_in_wlast(axi4frag_auto_in_wlast),
    .auto_in_bready(axi4frag_auto_in_bready),
    .auto_in_bvalid(axi4frag_auto_in_bvalid),
    .auto_in_bid(axi4frag_auto_in_bid),
    .auto_in_bresp(axi4frag_auto_in_bresp),
    .auto_in_buser(axi4frag_auto_in_buser),
    .auto_in_arready(axi4frag_auto_in_arready),
    .auto_in_arvalid(axi4frag_auto_in_arvalid),
    .auto_in_arid(axi4frag_auto_in_arid),
    .auto_in_araddr(axi4frag_auto_in_araddr),
    .auto_in_arlen(axi4frag_auto_in_arlen),
    .auto_in_arsize(axi4frag_auto_in_arsize),
    .auto_in_arburst(axi4frag_auto_in_arburst),
    .auto_in_aruser(axi4frag_auto_in_aruser),
    .auto_in_rready(axi4frag_auto_in_rready),
    .auto_in_rvalid(axi4frag_auto_in_rvalid),
    .auto_in_rid(axi4frag_auto_in_rid),
    .auto_in_rdata(axi4frag_auto_in_rdata),
    .auto_in_rresp(axi4frag_auto_in_rresp),
    .auto_in_ruser(axi4frag_auto_in_ruser),
    .auto_in_rlast(axi4frag_auto_in_rlast),
    .auto_out_awready(axi4frag_auto_out_awready),
    .auto_out_awvalid(axi4frag_auto_out_awvalid),
    .auto_out_awid(axi4frag_auto_out_awid),
    .auto_out_awaddr(axi4frag_auto_out_awaddr),
    .auto_out_awlen(axi4frag_auto_out_awlen),
    .auto_out_awsize(axi4frag_auto_out_awsize),
    .auto_out_awuser(axi4frag_auto_out_awuser),
    .auto_out_wready(axi4frag_auto_out_wready),
    .auto_out_wvalid(axi4frag_auto_out_wvalid),
    .auto_out_wdata(axi4frag_auto_out_wdata),
    .auto_out_wstrb(axi4frag_auto_out_wstrb),
    .auto_out_wlast(axi4frag_auto_out_wlast),
    .auto_out_bready(axi4frag_auto_out_bready),
    .auto_out_bvalid(axi4frag_auto_out_bvalid),
    .auto_out_bid(axi4frag_auto_out_bid),
    .auto_out_bresp(axi4frag_auto_out_bresp),
    .auto_out_buser(axi4frag_auto_out_buser),
    .auto_out_arready(axi4frag_auto_out_arready),
    .auto_out_arvalid(axi4frag_auto_out_arvalid),
    .auto_out_arid(axi4frag_auto_out_arid),
    .auto_out_araddr(axi4frag_auto_out_araddr),
    .auto_out_arlen(axi4frag_auto_out_arlen),
    .auto_out_arsize(axi4frag_auto_out_arsize),
    .auto_out_aruser(axi4frag_auto_out_aruser),
    .auto_out_rready(axi4frag_auto_out_rready),
    .auto_out_rvalid(axi4frag_auto_out_rvalid),
    .auto_out_rid(axi4frag_auto_out_rid),
    .auto_out_rdata(axi4frag_auto_out_rdata),
    .auto_out_rresp(axi4frag_auto_out_rresp),
    .auto_out_ruser(axi4frag_auto_out_ruser),
    .auto_out_rlast(axi4frag_auto_out_rlast)
  );
  dual_AXI4IdIndexer_2 axi4index_2 ( 
    .auto_in_awready(axi4index_2_auto_in_awready),
    .auto_in_awvalid(axi4index_2_auto_in_awvalid),
    .auto_in_awid(axi4index_2_auto_in_awid),
    .auto_in_awaddr(axi4index_2_auto_in_awaddr),
    .auto_in_awlen(axi4index_2_auto_in_awlen),
    .auto_in_awsize(axi4index_2_auto_in_awsize),
    .auto_in_awburst(axi4index_2_auto_in_awburst),
    .auto_in_wready(axi4index_2_auto_in_wready),
    .auto_in_wvalid(axi4index_2_auto_in_wvalid),
    .auto_in_wdata(axi4index_2_auto_in_wdata),
    .auto_in_wstrb(axi4index_2_auto_in_wstrb),
    .auto_in_wlast(axi4index_2_auto_in_wlast),
    .auto_in_bready(axi4index_2_auto_in_bready),
    .auto_in_bvalid(axi4index_2_auto_in_bvalid),
    .auto_in_bid(axi4index_2_auto_in_bid),
    .auto_in_bresp(axi4index_2_auto_in_bresp),
    .auto_in_arready(axi4index_2_auto_in_arready),
    .auto_in_arvalid(axi4index_2_auto_in_arvalid),
    .auto_in_arid(axi4index_2_auto_in_arid),
    .auto_in_araddr(axi4index_2_auto_in_araddr),
    .auto_in_arlen(axi4index_2_auto_in_arlen),
    .auto_in_arsize(axi4index_2_auto_in_arsize),
    .auto_in_arburst(axi4index_2_auto_in_arburst),
    .auto_in_rready(axi4index_2_auto_in_rready),
    .auto_in_rvalid(axi4index_2_auto_in_rvalid),
    .auto_in_rid(axi4index_2_auto_in_rid),
    .auto_in_rdata(axi4index_2_auto_in_rdata),
    .auto_in_rresp(axi4index_2_auto_in_rresp),
    .auto_in_rlast(axi4index_2_auto_in_rlast),
    .auto_out_awready(axi4index_2_auto_out_awready),
    .auto_out_awvalid(axi4index_2_auto_out_awvalid),
    .auto_out_awid(axi4index_2_auto_out_awid),
    .auto_out_awaddr(axi4index_2_auto_out_awaddr),
    .auto_out_awlen(axi4index_2_auto_out_awlen),
    .auto_out_awsize(axi4index_2_auto_out_awsize),
    .auto_out_awburst(axi4index_2_auto_out_awburst),
    .auto_out_awuser(axi4index_2_auto_out_awuser),
    .auto_out_wready(axi4index_2_auto_out_wready),
    .auto_out_wvalid(axi4index_2_auto_out_wvalid),
    .auto_out_wdata(axi4index_2_auto_out_wdata),
    .auto_out_wstrb(axi4index_2_auto_out_wstrb),
    .auto_out_wlast(axi4index_2_auto_out_wlast),
    .auto_out_bready(axi4index_2_auto_out_bready),
    .auto_out_bvalid(axi4index_2_auto_out_bvalid),
    .auto_out_bid(axi4index_2_auto_out_bid),
    .auto_out_bresp(axi4index_2_auto_out_bresp),
    .auto_out_buser(axi4index_2_auto_out_buser),
    .auto_out_arready(axi4index_2_auto_out_arready),
    .auto_out_arvalid(axi4index_2_auto_out_arvalid),
    .auto_out_arid(axi4index_2_auto_out_arid),
    .auto_out_araddr(axi4index_2_auto_out_araddr),
    .auto_out_arlen(axi4index_2_auto_out_arlen),
    .auto_out_arsize(axi4index_2_auto_out_arsize),
    .auto_out_arburst(axi4index_2_auto_out_arburst),
    .auto_out_aruser(axi4index_2_auto_out_aruser),
    .auto_out_rready(axi4index_2_auto_out_rready),
    .auto_out_rvalid(axi4index_2_auto_out_rvalid),
    .auto_out_rid(axi4index_2_auto_out_rid),
    .auto_out_rdata(axi4index_2_auto_out_rdata),
    .auto_out_rresp(axi4index_2_auto_out_rresp),
    .auto_out_ruser(axi4index_2_auto_out_ruser),
    .auto_out_rlast(axi4index_2_auto_out_rlast)
  );
  dual_TLError_2 err ( 
    .clock(err_clock),
    .reset(err_reset),
    .auto_in_a_ready(err_auto_in_a_ready),
    .auto_in_a_valid(err_auto_in_a_valid),
    .auto_in_a_bits_opcode(err_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(err_auto_in_a_bits_param),
    .auto_in_a_bits_size(err_auto_in_a_bits_size),
    .auto_in_a_bits_source(err_auto_in_a_bits_source),
    .auto_in_a_bits_address(err_auto_in_a_bits_address),
    .auto_in_a_bits_mask(err_auto_in_a_bits_mask),
    .auto_in_a_bits_corrupt(err_auto_in_a_bits_corrupt),
    .auto_in_c_ready(err_auto_in_c_ready),
    .auto_in_c_valid(err_auto_in_c_valid),
    .auto_in_c_bits_opcode(err_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(err_auto_in_c_bits_param),
    .auto_in_c_bits_size(err_auto_in_c_bits_size),
    .auto_in_c_bits_source(err_auto_in_c_bits_source),
    .auto_in_c_bits_address(err_auto_in_c_bits_address),
    .auto_in_c_bits_corrupt(err_auto_in_c_bits_corrupt),
    .auto_in_d_ready(err_auto_in_d_ready),
    .auto_in_d_valid(err_auto_in_d_valid),
    .auto_in_d_bits_opcode(err_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(err_auto_in_d_bits_param),
    .auto_in_d_bits_size(err_auto_in_d_bits_size),
    .auto_in_d_bits_source(err_auto_in_d_bits_source),
    .auto_in_d_bits_sink(err_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(err_auto_in_d_bits_denied),
    .auto_in_d_bits_data(err_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(err_auto_in_d_bits_corrupt),
    .auto_in_e_valid(err_auto_in_e_valid)
  );
  dual_TLAtomicAutomata atomics ( 
    .clock(atomics_clock),
    .reset(atomics_reset),
    .auto_in_a_ready(atomics_auto_in_a_ready),
    .auto_in_a_valid(atomics_auto_in_a_valid),
    .auto_in_a_bits_opcode(atomics_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(atomics_auto_in_a_bits_param),
    .auto_in_a_bits_size(atomics_auto_in_a_bits_size),
    .auto_in_a_bits_source(atomics_auto_in_a_bits_source),
    .auto_in_a_bits_address(atomics_auto_in_a_bits_address),
    .auto_in_a_bits_mask(atomics_auto_in_a_bits_mask),
    .auto_in_a_bits_data(atomics_auto_in_a_bits_data),
    .auto_in_c_ready(atomics_auto_in_c_ready),
    .auto_in_c_valid(atomics_auto_in_c_valid),
    .auto_in_c_bits_opcode(atomics_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(atomics_auto_in_c_bits_param),
    .auto_in_c_bits_size(atomics_auto_in_c_bits_size),
    .auto_in_c_bits_source(atomics_auto_in_c_bits_source),
    .auto_in_c_bits_address(atomics_auto_in_c_bits_address),
    .auto_in_c_bits_corrupt(atomics_auto_in_c_bits_corrupt),
    .auto_in_d_ready(atomics_auto_in_d_ready),
    .auto_in_d_valid(atomics_auto_in_d_valid),
    .auto_in_d_bits_opcode(atomics_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(atomics_auto_in_d_bits_param),
    .auto_in_d_bits_size(atomics_auto_in_d_bits_size),
    .auto_in_d_bits_source(atomics_auto_in_d_bits_source),
    .auto_in_d_bits_sink(atomics_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(atomics_auto_in_d_bits_denied),
    .auto_in_d_bits_data(atomics_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(atomics_auto_in_d_bits_corrupt),
    .auto_in_e_ready(atomics_auto_in_e_ready),
    .auto_in_e_valid(atomics_auto_in_e_valid),
    .auto_in_e_bits_sink(atomics_auto_in_e_bits_sink),
    .auto_out_a_ready(atomics_auto_out_a_ready),
    .auto_out_a_valid(atomics_auto_out_a_valid),
    .auto_out_a_bits_opcode(atomics_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(atomics_auto_out_a_bits_param),
    .auto_out_a_bits_size(atomics_auto_out_a_bits_size),
    .auto_out_a_bits_source(atomics_auto_out_a_bits_source),
    .auto_out_a_bits_address(atomics_auto_out_a_bits_address),
    .auto_out_a_bits_mask(atomics_auto_out_a_bits_mask),
    .auto_out_a_bits_data(atomics_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(atomics_auto_out_a_bits_corrupt),
    .auto_out_c_ready(atomics_auto_out_c_ready),
    .auto_out_c_valid(atomics_auto_out_c_valid),
    .auto_out_c_bits_opcode(atomics_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(atomics_auto_out_c_bits_param),
    .auto_out_c_bits_size(atomics_auto_out_c_bits_size),
    .auto_out_c_bits_source(atomics_auto_out_c_bits_source),
    .auto_out_c_bits_address(atomics_auto_out_c_bits_address),
    .auto_out_c_bits_corrupt(atomics_auto_out_c_bits_corrupt),
    .auto_out_d_ready(atomics_auto_out_d_ready),
    .auto_out_d_valid(atomics_auto_out_d_valid),
    .auto_out_d_bits_opcode(atomics_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(atomics_auto_out_d_bits_param),
    .auto_out_d_bits_size(atomics_auto_out_d_bits_size),
    .auto_out_d_bits_source(atomics_auto_out_d_bits_source),
    .auto_out_d_bits_sink(atomics_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(atomics_auto_out_d_bits_denied),
    .auto_out_d_bits_data(atomics_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(atomics_auto_out_d_bits_corrupt),
    .auto_out_e_ready(atomics_auto_out_e_ready),
    .auto_out_e_valid(atomics_auto_out_e_valid),
    .auto_out_e_bits_sink(atomics_auto_out_e_bits_sink)
  );
  dual_TLFIFOFixer_1 fixer_1 ( 
    .clock(fixer_1_clock),
    .reset(fixer_1_reset),
    .auto_in_a_ready(fixer_1_auto_in_a_ready),
    .auto_in_a_valid(fixer_1_auto_in_a_valid),
    .auto_in_a_bits_opcode(fixer_1_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(fixer_1_auto_in_a_bits_param),
    .auto_in_a_bits_size(fixer_1_auto_in_a_bits_size),
    .auto_in_a_bits_source(fixer_1_auto_in_a_bits_source),
    .auto_in_a_bits_address(fixer_1_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fixer_1_auto_in_a_bits_mask),
    .auto_in_a_bits_data(fixer_1_auto_in_a_bits_data),
    .auto_in_c_ready(fixer_1_auto_in_c_ready),
    .auto_in_c_valid(fixer_1_auto_in_c_valid),
    .auto_in_c_bits_opcode(fixer_1_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(fixer_1_auto_in_c_bits_param),
    .auto_in_c_bits_size(fixer_1_auto_in_c_bits_size),
    .auto_in_c_bits_source(fixer_1_auto_in_c_bits_source),
    .auto_in_c_bits_address(fixer_1_auto_in_c_bits_address),
    .auto_in_c_bits_corrupt(fixer_1_auto_in_c_bits_corrupt),
    .auto_in_d_ready(fixer_1_auto_in_d_ready),
    .auto_in_d_valid(fixer_1_auto_in_d_valid),
    .auto_in_d_bits_opcode(fixer_1_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(fixer_1_auto_in_d_bits_param),
    .auto_in_d_bits_size(fixer_1_auto_in_d_bits_size),
    .auto_in_d_bits_source(fixer_1_auto_in_d_bits_source),
    .auto_in_d_bits_sink(fixer_1_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(fixer_1_auto_in_d_bits_denied),
    .auto_in_d_bits_data(fixer_1_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(fixer_1_auto_in_d_bits_corrupt),
    .auto_in_e_ready(fixer_1_auto_in_e_ready),
    .auto_in_e_valid(fixer_1_auto_in_e_valid),
    .auto_in_e_bits_sink(fixer_1_auto_in_e_bits_sink),
    .auto_out_a_ready(fixer_1_auto_out_a_ready),
    .auto_out_a_valid(fixer_1_auto_out_a_valid),
    .auto_out_a_bits_opcode(fixer_1_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(fixer_1_auto_out_a_bits_param),
    .auto_out_a_bits_size(fixer_1_auto_out_a_bits_size),
    .auto_out_a_bits_source(fixer_1_auto_out_a_bits_source),
    .auto_out_a_bits_address(fixer_1_auto_out_a_bits_address),
    .auto_out_a_bits_mask(fixer_1_auto_out_a_bits_mask),
    .auto_out_a_bits_data(fixer_1_auto_out_a_bits_data),
    .auto_out_c_ready(fixer_1_auto_out_c_ready),
    .auto_out_c_valid(fixer_1_auto_out_c_valid),
    .auto_out_c_bits_opcode(fixer_1_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(fixer_1_auto_out_c_bits_param),
    .auto_out_c_bits_size(fixer_1_auto_out_c_bits_size),
    .auto_out_c_bits_source(fixer_1_auto_out_c_bits_source),
    .auto_out_c_bits_address(fixer_1_auto_out_c_bits_address),
    .auto_out_c_bits_corrupt(fixer_1_auto_out_c_bits_corrupt),
    .auto_out_d_ready(fixer_1_auto_out_d_ready),
    .auto_out_d_valid(fixer_1_auto_out_d_valid),
    .auto_out_d_bits_opcode(fixer_1_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(fixer_1_auto_out_d_bits_param),
    .auto_out_d_bits_size(fixer_1_auto_out_d_bits_size),
    .auto_out_d_bits_source(fixer_1_auto_out_d_bits_source),
    .auto_out_d_bits_sink(fixer_1_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(fixer_1_auto_out_d_bits_denied),
    .auto_out_d_bits_data(fixer_1_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(fixer_1_auto_out_d_bits_corrupt),
    .auto_out_e_ready(fixer_1_auto_out_e_ready),
    .auto_out_e_valid(fixer_1_auto_out_e_valid),
    .auto_out_e_bits_sink(fixer_1_auto_out_e_bits_sink)
  );
  dual_TLHintHandler hints ( 
    .clock(hints_clock),
    .reset(hints_reset),
    .auto_in_a_ready(hints_auto_in_a_ready),
    .auto_in_a_valid(hints_auto_in_a_valid),
    .auto_in_a_bits_opcode(hints_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(hints_auto_in_a_bits_param),
    .auto_in_a_bits_size(hints_auto_in_a_bits_size),
    .auto_in_a_bits_source(hints_auto_in_a_bits_source),
    .auto_in_a_bits_address(hints_auto_in_a_bits_address),
    .auto_in_a_bits_mask(hints_auto_in_a_bits_mask),
    .auto_in_a_bits_data(hints_auto_in_a_bits_data),
    .auto_in_c_ready(hints_auto_in_c_ready),
    .auto_in_c_valid(hints_auto_in_c_valid),
    .auto_in_c_bits_opcode(hints_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(hints_auto_in_c_bits_param),
    .auto_in_c_bits_size(hints_auto_in_c_bits_size),
    .auto_in_c_bits_source(hints_auto_in_c_bits_source),
    .auto_in_c_bits_address(hints_auto_in_c_bits_address),
    .auto_in_c_bits_corrupt(hints_auto_in_c_bits_corrupt),
    .auto_in_d_ready(hints_auto_in_d_ready),
    .auto_in_d_valid(hints_auto_in_d_valid),
    .auto_in_d_bits_opcode(hints_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(hints_auto_in_d_bits_param),
    .auto_in_d_bits_size(hints_auto_in_d_bits_size),
    .auto_in_d_bits_source(hints_auto_in_d_bits_source),
    .auto_in_d_bits_sink(hints_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(hints_auto_in_d_bits_denied),
    .auto_in_d_bits_data(hints_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(hints_auto_in_d_bits_corrupt),
    .auto_in_e_ready(hints_auto_in_e_ready),
    .auto_in_e_valid(hints_auto_in_e_valid),
    .auto_in_e_bits_sink(hints_auto_in_e_bits_sink),
    .auto_out_a_ready(hints_auto_out_a_ready),
    .auto_out_a_valid(hints_auto_out_a_valid),
    .auto_out_a_bits_opcode(hints_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(hints_auto_out_a_bits_param),
    .auto_out_a_bits_size(hints_auto_out_a_bits_size),
    .auto_out_a_bits_source(hints_auto_out_a_bits_source),
    .auto_out_a_bits_address(hints_auto_out_a_bits_address),
    .auto_out_a_bits_mask(hints_auto_out_a_bits_mask),
    .auto_out_a_bits_data(hints_auto_out_a_bits_data),
    .auto_out_c_ready(hints_auto_out_c_ready),
    .auto_out_c_valid(hints_auto_out_c_valid),
    .auto_out_c_bits_opcode(hints_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(hints_auto_out_c_bits_param),
    .auto_out_c_bits_size(hints_auto_out_c_bits_size),
    .auto_out_c_bits_source(hints_auto_out_c_bits_source),
    .auto_out_c_bits_address(hints_auto_out_c_bits_address),
    .auto_out_c_bits_corrupt(hints_auto_out_c_bits_corrupt),
    .auto_out_d_ready(hints_auto_out_d_ready),
    .auto_out_d_valid(hints_auto_out_d_valid),
    .auto_out_d_bits_opcode(hints_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(hints_auto_out_d_bits_param),
    .auto_out_d_bits_size(hints_auto_out_d_bits_size),
    .auto_out_d_bits_source(hints_auto_out_d_bits_source),
    .auto_out_d_bits_sink(hints_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(hints_auto_out_d_bits_denied),
    .auto_out_d_bits_data(hints_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(hints_auto_out_d_bits_corrupt),
    .auto_out_e_ready(hints_auto_out_e_ready),
    .auto_out_e_valid(hints_auto_out_e_valid),
    .auto_out_e_bits_sink(hints_auto_out_e_bits_sink)
  );
  dual_TLWidthWidget_1 widget_1 ( 
    .clock(widget_1_clock),
    .reset(widget_1_reset),
    .auto_in_a_ready(widget_1_auto_in_a_ready),
    .auto_in_a_valid(widget_1_auto_in_a_valid),
    .auto_in_a_bits_opcode(widget_1_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(widget_1_auto_in_a_bits_param),
    .auto_in_a_bits_size(widget_1_auto_in_a_bits_size),
    .auto_in_a_bits_source(widget_1_auto_in_a_bits_source),
    .auto_in_a_bits_address(widget_1_auto_in_a_bits_address),
    .auto_in_a_bits_mask(widget_1_auto_in_a_bits_mask),
    .auto_in_a_bits_data(widget_1_auto_in_a_bits_data),
    .auto_in_c_ready(widget_1_auto_in_c_ready),
    .auto_in_c_valid(widget_1_auto_in_c_valid),
    .auto_in_c_bits_opcode(widget_1_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(widget_1_auto_in_c_bits_param),
    .auto_in_c_bits_size(widget_1_auto_in_c_bits_size),
    .auto_in_c_bits_source(widget_1_auto_in_c_bits_source),
    .auto_in_c_bits_address(widget_1_auto_in_c_bits_address),
    .auto_in_c_bits_corrupt(widget_1_auto_in_c_bits_corrupt),
    .auto_in_d_ready(widget_1_auto_in_d_ready),
    .auto_in_d_valid(widget_1_auto_in_d_valid),
    .auto_in_d_bits_opcode(widget_1_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(widget_1_auto_in_d_bits_param),
    .auto_in_d_bits_size(widget_1_auto_in_d_bits_size),
    .auto_in_d_bits_source(widget_1_auto_in_d_bits_source),
    .auto_in_d_bits_sink(widget_1_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(widget_1_auto_in_d_bits_denied),
    .auto_in_d_bits_data(widget_1_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(widget_1_auto_in_d_bits_corrupt),
    .auto_in_e_ready(widget_1_auto_in_e_ready),
    .auto_in_e_valid(widget_1_auto_in_e_valid),
    .auto_in_e_bits_sink(widget_1_auto_in_e_bits_sink),
    .auto_out_a_ready(widget_1_auto_out_a_ready),
    .auto_out_a_valid(widget_1_auto_out_a_valid),
    .auto_out_a_bits_opcode(widget_1_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(widget_1_auto_out_a_bits_param),
    .auto_out_a_bits_size(widget_1_auto_out_a_bits_size),
    .auto_out_a_bits_source(widget_1_auto_out_a_bits_source),
    .auto_out_a_bits_address(widget_1_auto_out_a_bits_address),
    .auto_out_a_bits_mask(widget_1_auto_out_a_bits_mask),
    .auto_out_a_bits_data(widget_1_auto_out_a_bits_data),
    .auto_out_c_ready(widget_1_auto_out_c_ready),
    .auto_out_c_valid(widget_1_auto_out_c_valid),
    .auto_out_c_bits_opcode(widget_1_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(widget_1_auto_out_c_bits_param),
    .auto_out_c_bits_size(widget_1_auto_out_c_bits_size),
    .auto_out_c_bits_source(widget_1_auto_out_c_bits_source),
    .auto_out_c_bits_address(widget_1_auto_out_c_bits_address),
    .auto_out_c_bits_corrupt(widget_1_auto_out_c_bits_corrupt),
    .auto_out_d_ready(widget_1_auto_out_d_ready),
    .auto_out_d_valid(widget_1_auto_out_d_valid),
    .auto_out_d_bits_opcode(widget_1_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(widget_1_auto_out_d_bits_param),
    .auto_out_d_bits_size(widget_1_auto_out_d_bits_size),
    .auto_out_d_bits_source(widget_1_auto_out_d_bits_source),
    .auto_out_d_bits_sink(widget_1_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(widget_1_auto_out_d_bits_denied),
    .auto_out_d_bits_data(widget_1_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(widget_1_auto_out_d_bits_corrupt),
    .auto_out_e_ready(widget_1_auto_out_e_ready),
    .auto_out_e_valid(widget_1_auto_out_e_valid),
    .auto_out_e_bits_sink(widget_1_auto_out_e_bits_sink)
  );
  dual_TLWidthWidget_2 widget_2 ( 
    .clock(widget_2_clock),
    .reset(widget_2_reset),
    .auto_in_a_ready(widget_2_auto_in_a_ready),
    .auto_in_a_valid(widget_2_auto_in_a_valid),
    .auto_in_a_bits_opcode(widget_2_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(widget_2_auto_in_a_bits_param),
    .auto_in_a_bits_size(widget_2_auto_in_a_bits_size),
    .auto_in_a_bits_source(widget_2_auto_in_a_bits_source),
    .auto_in_a_bits_address(widget_2_auto_in_a_bits_address),
    .auto_in_a_bits_mask(widget_2_auto_in_a_bits_mask),
    .auto_in_a_bits_corrupt(widget_2_auto_in_a_bits_corrupt),
    .auto_in_c_ready(widget_2_auto_in_c_ready),
    .auto_in_c_valid(widget_2_auto_in_c_valid),
    .auto_in_c_bits_opcode(widget_2_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(widget_2_auto_in_c_bits_param),
    .auto_in_c_bits_size(widget_2_auto_in_c_bits_size),
    .auto_in_c_bits_source(widget_2_auto_in_c_bits_source),
    .auto_in_c_bits_address(widget_2_auto_in_c_bits_address),
    .auto_in_c_bits_corrupt(widget_2_auto_in_c_bits_corrupt),
    .auto_in_d_ready(widget_2_auto_in_d_ready),
    .auto_in_d_valid(widget_2_auto_in_d_valid),
    .auto_in_d_bits_opcode(widget_2_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(widget_2_auto_in_d_bits_param),
    .auto_in_d_bits_size(widget_2_auto_in_d_bits_size),
    .auto_in_d_bits_source(widget_2_auto_in_d_bits_source),
    .auto_in_d_bits_sink(widget_2_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(widget_2_auto_in_d_bits_denied),
    .auto_in_d_bits_data(widget_2_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(widget_2_auto_in_d_bits_corrupt),
    .auto_in_e_valid(widget_2_auto_in_e_valid),
    .auto_out_a_ready(widget_2_auto_out_a_ready),
    .auto_out_a_valid(widget_2_auto_out_a_valid),
    .auto_out_a_bits_opcode(widget_2_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(widget_2_auto_out_a_bits_param),
    .auto_out_a_bits_size(widget_2_auto_out_a_bits_size),
    .auto_out_a_bits_source(widget_2_auto_out_a_bits_source),
    .auto_out_a_bits_address(widget_2_auto_out_a_bits_address),
    .auto_out_a_bits_mask(widget_2_auto_out_a_bits_mask),
    .auto_out_a_bits_corrupt(widget_2_auto_out_a_bits_corrupt),
    .auto_out_c_ready(widget_2_auto_out_c_ready),
    .auto_out_c_valid(widget_2_auto_out_c_valid),
    .auto_out_c_bits_opcode(widget_2_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(widget_2_auto_out_c_bits_param),
    .auto_out_c_bits_size(widget_2_auto_out_c_bits_size),
    .auto_out_c_bits_source(widget_2_auto_out_c_bits_source),
    .auto_out_c_bits_address(widget_2_auto_out_c_bits_address),
    .auto_out_c_bits_corrupt(widget_2_auto_out_c_bits_corrupt),
    .auto_out_d_ready(widget_2_auto_out_d_ready),
    .auto_out_d_valid(widget_2_auto_out_d_valid),
    .auto_out_d_bits_opcode(widget_2_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(widget_2_auto_out_d_bits_param),
    .auto_out_d_bits_size(widget_2_auto_out_d_bits_size),
    .auto_out_d_bits_source(widget_2_auto_out_d_bits_source),
    .auto_out_d_bits_sink(widget_2_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(widget_2_auto_out_d_bits_denied),
    .auto_out_d_bits_data(widget_2_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(widget_2_auto_out_d_bits_corrupt),
    .auto_out_e_valid(widget_2_auto_out_e_valid)
  );
  assign fpga_io_c2b_clk = chiplink_auto_io_out_c2b_clk; 
  assign fpga_io_c2b_rst = chiplink_auto_io_out_c2b_rst; 
  assign fpga_io_c2b_send = chiplink_auto_io_out_c2b_send; 
  assign fpga_io_c2b_data = chiplink_auto_io_out_c2b_data; 
  assign mem_axi4_0_awvalid = axi4yank_auto_out_awvalid; 
  assign mem_axi4_0_awid = axi4yank_auto_out_awid; 
  assign mem_axi4_0_awaddr = axi4yank_auto_out_awaddr; 
  assign mem_axi4_0_awlen = axi4yank_auto_out_awlen; 
  assign mem_axi4_0_awsize = axi4yank_auto_out_awsize; 
  assign mem_axi4_0_awburst = axi4yank_auto_out_awburst; 
  assign mem_axi4_0_awlock = axi4yank_auto_out_awlock; 
  assign mem_axi4_0_awcache = axi4yank_auto_out_awcache; 
  assign mem_axi4_0_awprot = axi4yank_auto_out_awprot; 
  assign mem_axi4_0_awqos = axi4yank_auto_out_awqos; 
  assign mem_axi4_0_awinstret = axi4yank_auto_out_awinstret; 
  assign mem_axi4_0_wvalid = axi4yank_auto_out_wvalid; 
  assign mem_axi4_0_wdata = axi4yank_auto_out_wdata; 
  assign mem_axi4_0_wstrb = axi4yank_auto_out_wstrb; 
  assign mem_axi4_0_wlast = axi4yank_auto_out_wlast; 
  assign mem_axi4_0_bready = axi4yank_auto_out_bready; 
  assign mem_axi4_0_arvalid = axi4yank_auto_out_arvalid; 
  assign mem_axi4_0_arid = axi4yank_auto_out_arid; 
  assign mem_axi4_0_araddr = axi4yank_auto_out_araddr; 
  assign mem_axi4_0_arlen = axi4yank_auto_out_arlen; 
  assign mem_axi4_0_arsize = axi4yank_auto_out_arsize; 
  assign mem_axi4_0_arburst = axi4yank_auto_out_arburst; 
  assign mem_axi4_0_arlock = axi4yank_auto_out_arlock; 
  assign mem_axi4_0_arcache = axi4yank_auto_out_arcache; 
  assign mem_axi4_0_arprot = axi4yank_auto_out_arprot; 
  assign mem_axi4_0_arqos = axi4yank_auto_out_arqos; 
  assign mem_axi4_0_arinstret = axi4yank_auto_out_arinstret; 
  assign mem_axi4_0_rready = axi4yank_auto_out_rready; 
  assign mmio_axi4_0_awvalid = axi4buf_auto_out_awvalid; 
  assign mmio_axi4_0_awid = axi4buf_auto_out_awid; 
  assign mmio_axi4_0_awaddr = axi4buf_auto_out_awaddr; 
  assign mmio_axi4_0_awlen = axi4buf_auto_out_awlen; 
  assign mmio_axi4_0_awsize = axi4buf_auto_out_awsize; 
  assign mmio_axi4_0_awburst = axi4buf_auto_out_awburst; 
  assign mmio_axi4_0_awlock = axi4buf_auto_out_awlock; 
  assign mmio_axi4_0_awcache = axi4buf_auto_out_awcache; 
  assign mmio_axi4_0_awprot = axi4buf_auto_out_awprot; 
  assign mmio_axi4_0_awqos = axi4buf_auto_out_awqos; 
  assign mmio_axi4_0_awinstret = axi4buf_auto_out_awinstret; 
  assign mmio_axi4_0_wvalid = axi4buf_auto_out_wvalid; 
  assign mmio_axi4_0_wdata = axi4buf_auto_out_wdata; 
  assign mmio_axi4_0_wstrb = axi4buf_auto_out_wstrb; 
  assign mmio_axi4_0_wlast = axi4buf_auto_out_wlast; 
  assign mmio_axi4_0_bready = axi4buf_auto_out_bready; 
  assign mmio_axi4_0_arvalid = axi4buf_auto_out_arvalid; 
  assign mmio_axi4_0_arid = axi4buf_auto_out_arid; 
  assign mmio_axi4_0_araddr = axi4buf_auto_out_araddr; 
  assign mmio_axi4_0_arlen = axi4buf_auto_out_arlen; 
  assign mmio_axi4_0_arsize = axi4buf_auto_out_arsize; 
  assign mmio_axi4_0_arburst = axi4buf_auto_out_arburst; 
  assign mmio_axi4_0_arlock = axi4buf_auto_out_arlock; 
  assign mmio_axi4_0_arcache = axi4buf_auto_out_arcache; 
  assign mmio_axi4_0_arprot = axi4buf_auto_out_arprot; 
  assign mmio_axi4_0_arqos = axi4buf_auto_out_arqos; 
  assign mmio_axi4_0_arinstret = axi4buf_auto_out_arinstret; 
  assign mmio_axi4_0_rready = axi4buf_auto_out_rready; 
  assign l2_frontend_bus_axi4_0_awready = axi4index_2_auto_in_awready; 
  assign l2_frontend_bus_axi4_0_wready = axi4index_2_auto_in_wready; 
  assign l2_frontend_bus_axi4_0_bvalid = axi4index_2_auto_in_bvalid; 
  assign l2_frontend_bus_axi4_0_bid = axi4index_2_auto_in_bid; 
  assign l2_frontend_bus_axi4_0_bresp = axi4index_2_auto_in_bresp; 
  assign l2_frontend_bus_axi4_0_arready = axi4index_2_auto_in_arready; 
  assign l2_frontend_bus_axi4_0_rvalid = axi4index_2_auto_in_rvalid; 
  assign l2_frontend_bus_axi4_0_rid = axi4index_2_auto_in_rid; 
  assign l2_frontend_bus_axi4_0_rdata = axi4index_2_auto_in_rdata; 
  assign l2_frontend_bus_axi4_0_rresp = axi4index_2_auto_in_rresp; 
  assign l2_frontend_bus_axi4_0_rlast = axi4index_2_auto_in_rlast; 
  assign xbar_clock = clock; 
  assign xbar_reset = reset; 
  assign xbar_auto_in_a_valid = atomics_auto_out_a_valid; 
  assign xbar_auto_in_a_bits_opcode = atomics_auto_out_a_bits_opcode; 
  assign xbar_auto_in_a_bits_param = atomics_auto_out_a_bits_param; 
  assign xbar_auto_in_a_bits_size = atomics_auto_out_a_bits_size; 
  assign xbar_auto_in_a_bits_source = atomics_auto_out_a_bits_source; 
  assign xbar_auto_in_a_bits_address = atomics_auto_out_a_bits_address; 
  assign xbar_auto_in_a_bits_mask = atomics_auto_out_a_bits_mask; 
  assign xbar_auto_in_a_bits_data = atomics_auto_out_a_bits_data; 
  assign xbar_auto_in_a_bits_corrupt = atomics_auto_out_a_bits_corrupt; 
  assign xbar_auto_in_c_valid = atomics_auto_out_c_valid; 
  assign xbar_auto_in_c_bits_opcode = atomics_auto_out_c_bits_opcode; 
  assign xbar_auto_in_c_bits_param = atomics_auto_out_c_bits_param; 
  assign xbar_auto_in_c_bits_size = atomics_auto_out_c_bits_size; 
  assign xbar_auto_in_c_bits_source = atomics_auto_out_c_bits_source; 
  assign xbar_auto_in_c_bits_address = atomics_auto_out_c_bits_address; 
  assign xbar_auto_in_c_bits_corrupt = atomics_auto_out_c_bits_corrupt; 
  assign xbar_auto_in_d_ready = atomics_auto_out_d_ready; 
  assign xbar_auto_in_e_valid = atomics_auto_out_e_valid; 
  assign xbar_auto_in_e_bits_sink = atomics_auto_out_e_bits_sink; 
  assign xbar_auto_out_2_a_ready = widget_2_auto_in_a_ready; 
  assign xbar_auto_out_2_c_ready = widget_2_auto_in_c_ready; 
  assign xbar_auto_out_2_d_valid = widget_2_auto_in_d_valid; 
  assign xbar_auto_out_2_d_bits_opcode = widget_2_auto_in_d_bits_opcode; 
  assign xbar_auto_out_2_d_bits_param = widget_2_auto_in_d_bits_param; 
  assign xbar_auto_out_2_d_bits_size = widget_2_auto_in_d_bits_size; 
  assign xbar_auto_out_2_d_bits_source = widget_2_auto_in_d_bits_source; 
  assign xbar_auto_out_2_d_bits_sink = widget_2_auto_in_d_bits_sink; 
  assign xbar_auto_out_2_d_bits_denied = widget_2_auto_in_d_bits_denied; 
  assign xbar_auto_out_2_d_bits_data = widget_2_auto_in_d_bits_data; 
  assign xbar_auto_out_2_d_bits_corrupt = widget_2_auto_in_d_bits_corrupt; 
  assign xbar_auto_out_1_a_ready = tl2axi4_1_auto_in_a_ready; 
  assign xbar_auto_out_1_d_valid = tl2axi4_1_auto_in_d_valid; 
  assign xbar_auto_out_1_d_bits_opcode = tl2axi4_1_auto_in_d_bits_opcode; 
  assign xbar_auto_out_1_d_bits_size = tl2axi4_1_auto_in_d_bits_size; 
  assign xbar_auto_out_1_d_bits_source = tl2axi4_1_auto_in_d_bits_source; 
  assign xbar_auto_out_1_d_bits_denied = tl2axi4_1_auto_in_d_bits_denied; 
  assign xbar_auto_out_1_d_bits_data = tl2axi4_1_auto_in_d_bits_data; 
  assign xbar_auto_out_1_d_bits_corrupt = tl2axi4_1_auto_in_d_bits_corrupt; 
  assign xbar_auto_out_0_a_ready = tl2axi4_auto_in_a_ready; 
  assign xbar_auto_out_0_d_valid = tl2axi4_auto_in_d_valid; 
  assign xbar_auto_out_0_d_bits_opcode = tl2axi4_auto_in_d_bits_opcode; 
  assign xbar_auto_out_0_d_bits_size = tl2axi4_auto_in_d_bits_size; 
  assign xbar_auto_out_0_d_bits_source = tl2axi4_auto_in_d_bits_source; 
  assign xbar_auto_out_0_d_bits_denied = tl2axi4_auto_in_d_bits_denied; 
  assign xbar_auto_out_0_d_bits_data = tl2axi4_auto_in_d_bits_data; 
  assign xbar_auto_out_0_d_bits_corrupt = tl2axi4_auto_in_d_bits_corrupt; 
  assign xbar_1_clock = clock; 
  assign xbar_1_reset = reset; 
  assign xbar_1_auto_in_a_valid = fixer_auto_out_a_valid; 
  assign xbar_1_auto_in_a_bits_opcode = fixer_auto_out_a_bits_opcode; 
  assign xbar_1_auto_in_a_bits_param = fixer_auto_out_a_bits_param; 
  assign xbar_1_auto_in_a_bits_size = fixer_auto_out_a_bits_size; 
  assign xbar_1_auto_in_a_bits_source = fixer_auto_out_a_bits_source; 
  assign xbar_1_auto_in_a_bits_address = fixer_auto_out_a_bits_address; 
  assign xbar_1_auto_in_a_bits_mask = fixer_auto_out_a_bits_mask; 
  assign xbar_1_auto_in_a_bits_data = fixer_auto_out_a_bits_data; 
  assign xbar_1_auto_in_a_bits_corrupt = fixer_auto_out_a_bits_corrupt; 
  assign xbar_1_auto_in_d_ready = fixer_auto_out_d_ready; 
  assign xbar_1_auto_out_1_a_ready = ferr_auto_in_a_ready; 
  assign xbar_1_auto_out_1_d_valid = ferr_auto_in_d_valid; 
  assign xbar_1_auto_out_1_d_bits_opcode = ferr_auto_in_d_bits_opcode; 
  assign xbar_1_auto_out_1_d_bits_param = ferr_auto_in_d_bits_param; 
  assign xbar_1_auto_out_1_d_bits_size = ferr_auto_in_d_bits_size; 
  assign xbar_1_auto_out_1_d_bits_source = ferr_auto_in_d_bits_source; 
  assign xbar_1_auto_out_1_d_bits_sink = ferr_auto_in_d_bits_sink; 
  assign xbar_1_auto_out_1_d_bits_denied = ferr_auto_in_d_bits_denied; 
  assign xbar_1_auto_out_1_d_bits_data = ferr_auto_in_d_bits_data; 
  assign xbar_1_auto_out_1_d_bits_corrupt = ferr_auto_in_d_bits_corrupt; 
  assign xbar_1_auto_out_0_a_ready = chiplink_auto_sbypass_node_in_in_a_ready; 
  assign xbar_1_auto_out_0_d_valid = chiplink_auto_sbypass_node_in_in_d_valid; 
  assign xbar_1_auto_out_0_d_bits_opcode = chiplink_auto_sbypass_node_in_in_d_bits_opcode; 
  assign xbar_1_auto_out_0_d_bits_param = chiplink_auto_sbypass_node_in_in_d_bits_param; 
  assign xbar_1_auto_out_0_d_bits_size = chiplink_auto_sbypass_node_in_in_d_bits_size; 
  assign xbar_1_auto_out_0_d_bits_source = chiplink_auto_sbypass_node_in_in_d_bits_source; 
  assign xbar_1_auto_out_0_d_bits_sink = chiplink_auto_sbypass_node_in_in_d_bits_sink; 
  assign xbar_1_auto_out_0_d_bits_denied = chiplink_auto_sbypass_node_in_in_d_bits_denied; 
  assign xbar_1_auto_out_0_d_bits_data = chiplink_auto_sbypass_node_in_in_d_bits_data; 
  assign xbar_1_auto_out_0_d_bits_corrupt = chiplink_auto_sbypass_node_in_in_d_bits_corrupt; 
  assign ferr_clock = clock; 
  assign ferr_reset = reset; 
  assign ferr_auto_in_a_valid = xbar_1_auto_out_1_a_valid; 
  assign ferr_auto_in_a_bits_opcode = xbar_1_auto_out_1_a_bits_opcode; 
  assign ferr_auto_in_a_bits_param = xbar_1_auto_out_1_a_bits_param; 
  assign ferr_auto_in_a_bits_size = xbar_1_auto_out_1_a_bits_size; 
  assign ferr_auto_in_a_bits_source = xbar_1_auto_out_1_a_bits_source; 
  assign ferr_auto_in_a_bits_address = xbar_1_auto_out_1_a_bits_address; 
  assign ferr_auto_in_a_bits_mask = xbar_1_auto_out_1_a_bits_mask; 
  assign ferr_auto_in_a_bits_corrupt = xbar_1_auto_out_1_a_bits_corrupt; 
  assign ferr_auto_in_d_ready = xbar_1_auto_out_1_d_ready; 
  assign chiplink_clock = clock; 
  assign chiplink_reset = reset; 
  assign chiplink_auto_mbypass_out_a_ready = widget_1_auto_in_a_ready; 
  assign chiplink_auto_mbypass_out_c_ready = widget_1_auto_in_c_ready; 
  assign chiplink_auto_mbypass_out_d_valid = widget_1_auto_in_d_valid; 
  assign chiplink_auto_mbypass_out_d_bits_opcode = widget_1_auto_in_d_bits_opcode; 
  assign chiplink_auto_mbypass_out_d_bits_param = widget_1_auto_in_d_bits_param; 
  assign chiplink_auto_mbypass_out_d_bits_size = widget_1_auto_in_d_bits_size; 
  assign chiplink_auto_mbypass_out_d_bits_source = widget_1_auto_in_d_bits_source; 
  assign chiplink_auto_mbypass_out_d_bits_sink = widget_1_auto_in_d_bits_sink; 
  assign chiplink_auto_mbypass_out_d_bits_denied = widget_1_auto_in_d_bits_denied; 
  assign chiplink_auto_mbypass_out_d_bits_data = widget_1_auto_in_d_bits_data; 
  assign chiplink_auto_mbypass_out_d_bits_corrupt = widget_1_auto_in_d_bits_corrupt; 
  assign chiplink_auto_mbypass_out_e_ready = widget_1_auto_in_e_ready; 
  assign chiplink_auto_sbypass_node_in_in_a_valid = xbar_1_auto_out_0_a_valid; 
  assign chiplink_auto_sbypass_node_in_in_a_bits_opcode = xbar_1_auto_out_0_a_bits_opcode; 
  assign chiplink_auto_sbypass_node_in_in_a_bits_param = xbar_1_auto_out_0_a_bits_param; 
  assign chiplink_auto_sbypass_node_in_in_a_bits_size = xbar_1_auto_out_0_a_bits_size; 
  assign chiplink_auto_sbypass_node_in_in_a_bits_source = xbar_1_auto_out_0_a_bits_source; 
  assign chiplink_auto_sbypass_node_in_in_a_bits_address = xbar_1_auto_out_0_a_bits_address; 
  assign chiplink_auto_sbypass_node_in_in_a_bits_mask = xbar_1_auto_out_0_a_bits_mask; 
  assign chiplink_auto_sbypass_node_in_in_a_bits_data = xbar_1_auto_out_0_a_bits_data; 
  assign chiplink_auto_sbypass_node_in_in_a_bits_corrupt = xbar_1_auto_out_0_a_bits_corrupt; 
  assign chiplink_auto_sbypass_node_in_in_d_ready = xbar_1_auto_out_0_d_ready; 
  assign chiplink_auto_io_out_b2c_clk = fpga_io_b2c_clk; 
  assign chiplink_auto_io_out_b2c_rst = fpga_io_b2c_rst; 
  assign chiplink_auto_io_out_b2c_send = fpga_io_b2c_send; 
  assign chiplink_auto_io_out_b2c_data = fpga_io_b2c_data; 
  assign axi4yank_clock = clock; 
  assign axi4yank_reset = reset; 
  assign axi4yank_auto_in_awvalid = axi4index_auto_out_awvalid; 
  assign axi4yank_auto_in_awid = axi4index_auto_out_awid; 
  assign axi4yank_auto_in_awaddr = axi4index_auto_out_awaddr; 
  assign axi4yank_auto_in_awlen = axi4index_auto_out_awlen; 
  assign axi4yank_auto_in_awsize = axi4index_auto_out_awsize; 
  assign axi4yank_auto_in_awburst = axi4index_auto_out_awburst; 
  assign axi4yank_auto_in_awlock = axi4index_auto_out_awlock; 
  assign axi4yank_auto_in_awcache = axi4index_auto_out_awcache; 
  assign axi4yank_auto_in_awprot = axi4index_auto_out_awprot; 
  assign axi4yank_auto_in_awqos = axi4index_auto_out_awqos; 
  assign axi4yank_auto_in_awuser = axi4index_auto_out_awuser; 
  assign axi4yank_auto_in_awinstret = axi4index_auto_out_awinstret; 
  assign axi4yank_auto_in_wvalid = axi4index_auto_out_wvalid; 
  assign axi4yank_auto_in_wdata = axi4index_auto_out_wdata; 
  assign axi4yank_auto_in_wstrb = axi4index_auto_out_wstrb; 
  assign axi4yank_auto_in_wlast = axi4index_auto_out_wlast; 
  assign axi4yank_auto_in_bready = axi4index_auto_out_bready; 
  assign axi4yank_auto_in_arvalid = axi4index_auto_out_arvalid; 
  assign axi4yank_auto_in_arid = axi4index_auto_out_arid; 
  assign axi4yank_auto_in_araddr = axi4index_auto_out_araddr; 
  assign axi4yank_auto_in_arlen = axi4index_auto_out_arlen; 
  assign axi4yank_auto_in_arsize = axi4index_auto_out_arsize; 
  assign axi4yank_auto_in_arburst = axi4index_auto_out_arburst; 
  assign axi4yank_auto_in_arlock = axi4index_auto_out_arlock; 
  assign axi4yank_auto_in_arcache = axi4index_auto_out_arcache; 
  assign axi4yank_auto_in_arprot = axi4index_auto_out_arprot; 
  assign axi4yank_auto_in_arqos = axi4index_auto_out_arqos; 
  assign axi4yank_auto_in_aruser = axi4index_auto_out_aruser; 
  assign axi4yank_auto_in_arinstret = axi4index_auto_out_arinstret; 
  assign axi4yank_auto_in_rready = axi4index_auto_out_rready; 
  assign axi4yank_auto_out_awready = mem_axi4_0_awready; 
  assign axi4yank_auto_out_wready = mem_axi4_0_wready; 
  assign axi4yank_auto_out_bvalid = mem_axi4_0_bvalid; 
  assign axi4yank_auto_out_bid = mem_axi4_0_bid; 
  assign axi4yank_auto_out_bresp = mem_axi4_0_bresp; 
  assign axi4yank_auto_out_arready = mem_axi4_0_arready; 
  assign axi4yank_auto_out_rvalid = mem_axi4_0_rvalid; 
  assign axi4yank_auto_out_rid = mem_axi4_0_rid; 
  assign axi4yank_auto_out_rdata = mem_axi4_0_rdata; 
  assign axi4yank_auto_out_rresp = mem_axi4_0_rresp; 
  assign axi4yank_auto_out_rlast = mem_axi4_0_rlast; 
  assign axi4index_auto_in_awvalid = tl2axi4_auto_out_awvalid; 
  assign axi4index_auto_in_awid = tl2axi4_auto_out_awid; 
  assign axi4index_auto_in_awaddr = tl2axi4_auto_out_awaddr; 
  assign axi4index_auto_in_awlen = tl2axi4_auto_out_awlen; 
  assign axi4index_auto_in_awsize = tl2axi4_auto_out_awsize; 
  assign axi4index_auto_in_awburst = tl2axi4_auto_out_awburst; 
  assign axi4index_auto_in_awlock = tl2axi4_auto_out_awlock; 
  assign axi4index_auto_in_awcache = tl2axi4_auto_out_awcache; 
  assign axi4index_auto_in_awprot = tl2axi4_auto_out_awprot; 
  assign axi4index_auto_in_awqos = tl2axi4_auto_out_awqos; 
  assign axi4index_auto_in_awuser = tl2axi4_auto_out_awuser; 
  assign axi4index_auto_in_awinstret = tl2axi4_auto_out_awinstret; 
  assign axi4index_auto_in_wvalid = tl2axi4_auto_out_wvalid; 
  assign axi4index_auto_in_wdata = tl2axi4_auto_out_wdata; 
  assign axi4index_auto_in_wstrb = tl2axi4_auto_out_wstrb; 
  assign axi4index_auto_in_wlast = tl2axi4_auto_out_wlast; 
  assign axi4index_auto_in_bready = tl2axi4_auto_out_bready; 
  assign axi4index_auto_in_arvalid = tl2axi4_auto_out_arvalid; 
  assign axi4index_auto_in_arid = tl2axi4_auto_out_arid; 
  assign axi4index_auto_in_araddr = tl2axi4_auto_out_araddr; 
  assign axi4index_auto_in_arlen = tl2axi4_auto_out_arlen; 
  assign axi4index_auto_in_arsize = tl2axi4_auto_out_arsize; 
  assign axi4index_auto_in_arburst = tl2axi4_auto_out_arburst; 
  assign axi4index_auto_in_arlock = tl2axi4_auto_out_arlock; 
  assign axi4index_auto_in_arcache = tl2axi4_auto_out_arcache; 
  assign axi4index_auto_in_arprot = tl2axi4_auto_out_arprot; 
  assign axi4index_auto_in_arqos = tl2axi4_auto_out_arqos; 
  assign axi4index_auto_in_aruser = tl2axi4_auto_out_aruser; 
  assign axi4index_auto_in_arinstret = tl2axi4_auto_out_arinstret; 
  assign axi4index_auto_in_rready = tl2axi4_auto_out_rready; 
  assign axi4index_auto_out_awready = axi4yank_auto_in_awready; 
  assign axi4index_auto_out_wready = axi4yank_auto_in_wready; 
  assign axi4index_auto_out_bvalid = axi4yank_auto_in_bvalid; 
  assign axi4index_auto_out_bid = axi4yank_auto_in_bid; 
  assign axi4index_auto_out_bresp = axi4yank_auto_in_bresp; 
  assign axi4index_auto_out_buser = axi4yank_auto_in_buser; 
  assign axi4index_auto_out_arready = axi4yank_auto_in_arready; 
  assign axi4index_auto_out_rvalid = axi4yank_auto_in_rvalid; 
  assign axi4index_auto_out_rid = axi4yank_auto_in_rid; 
  assign axi4index_auto_out_rdata = axi4yank_auto_in_rdata; 
  assign axi4index_auto_out_rresp = axi4yank_auto_in_rresp; 
  assign axi4index_auto_out_ruser = axi4yank_auto_in_ruser; 
  assign axi4index_auto_out_rlast = axi4yank_auto_in_rlast; 
  assign tl2axi4_clock = clock; 
  assign tl2axi4_reset = reset; 
  assign tl2axi4_auto_in_a_valid = xbar_auto_out_0_a_valid; 
  assign tl2axi4_auto_in_a_bits_opcode = xbar_auto_out_0_a_bits_opcode; 
  assign tl2axi4_auto_in_a_bits_param = xbar_auto_out_0_a_bits_param; 
  assign tl2axi4_auto_in_a_bits_size = xbar_auto_out_0_a_bits_size; 
  assign tl2axi4_auto_in_a_bits_source = xbar_auto_out_0_a_bits_source; 
  assign tl2axi4_auto_in_a_bits_address = xbar_auto_out_0_a_bits_address; 
  assign tl2axi4_auto_in_a_bits_mask = xbar_auto_out_0_a_bits_mask; 
  assign tl2axi4_auto_in_a_bits_data = xbar_auto_out_0_a_bits_data; 
  assign tl2axi4_auto_in_a_bits_corrupt = xbar_auto_out_0_a_bits_corrupt; 
  assign tl2axi4_auto_in_d_ready = xbar_auto_out_0_d_ready; 
  assign tl2axi4_auto_out_awready = axi4index_auto_in_awready; 
  assign tl2axi4_auto_out_wready = axi4index_auto_in_wready; 
  assign tl2axi4_auto_out_bvalid = axi4index_auto_in_bvalid; 
  assign tl2axi4_auto_out_bid = axi4index_auto_in_bid; 
  assign tl2axi4_auto_out_bresp = axi4index_auto_in_bresp; 
  assign tl2axi4_auto_out_buser = axi4index_auto_in_buser; 
  assign tl2axi4_auto_out_arready = axi4index_auto_in_arready; 
  assign tl2axi4_auto_out_rvalid = axi4index_auto_in_rvalid; 
  assign tl2axi4_auto_out_rid = axi4index_auto_in_rid; 
  assign tl2axi4_auto_out_rdata = axi4index_auto_in_rdata; 
  assign tl2axi4_auto_out_rresp = axi4index_auto_in_rresp; 
  assign tl2axi4_auto_out_ruser = axi4index_auto_in_ruser; 
  assign tl2axi4_auto_out_rlast = axi4index_auto_in_rlast; 
  assign axi4buf_clock = clock; 
  assign axi4buf_reset = reset; 
  assign axi4buf_auto_in_awvalid = axi4yank_1_auto_out_awvalid; 
  assign axi4buf_auto_in_awaddr = axi4yank_1_auto_out_awaddr; 
  assign axi4buf_auto_in_awlen = axi4yank_1_auto_out_awlen; 
  assign axi4buf_auto_in_awsize = axi4yank_1_auto_out_awsize; 
  assign axi4buf_auto_in_awburst = axi4yank_1_auto_out_awburst; 
  assign axi4buf_auto_in_awlock = axi4yank_1_auto_out_awlock; 
  assign axi4buf_auto_in_awcache = axi4yank_1_auto_out_awcache; 
  assign axi4buf_auto_in_awprot = axi4yank_1_auto_out_awprot; 
  assign axi4buf_auto_in_awqos = axi4yank_1_auto_out_awqos; 
  assign axi4buf_auto_in_awinstret = axi4yank_1_auto_out_awinstret; 
  assign axi4buf_auto_in_wvalid = axi4yank_1_auto_out_wvalid; 
  assign axi4buf_auto_in_wdata = axi4yank_1_auto_out_wdata; 
  assign axi4buf_auto_in_wstrb = axi4yank_1_auto_out_wstrb; 
  assign axi4buf_auto_in_wlast = axi4yank_1_auto_out_wlast; 
  assign axi4buf_auto_in_bready = axi4yank_1_auto_out_bready; 
  assign axi4buf_auto_in_arvalid = axi4yank_1_auto_out_arvalid; 
  assign axi4buf_auto_in_araddr = axi4yank_1_auto_out_araddr; 
  assign axi4buf_auto_in_arlen = axi4yank_1_auto_out_arlen; 
  assign axi4buf_auto_in_arsize = axi4yank_1_auto_out_arsize; 
  assign axi4buf_auto_in_arburst = axi4yank_1_auto_out_arburst; 
  assign axi4buf_auto_in_arlock = axi4yank_1_auto_out_arlock; 
  assign axi4buf_auto_in_arcache = axi4yank_1_auto_out_arcache; 
  assign axi4buf_auto_in_arprot = axi4yank_1_auto_out_arprot; 
  assign axi4buf_auto_in_arqos = axi4yank_1_auto_out_arqos; 
  assign axi4buf_auto_in_arinstret = axi4yank_1_auto_out_arinstret; 
  assign axi4buf_auto_in_rready = axi4yank_1_auto_out_rready; 
  assign axi4buf_auto_out_awready = mmio_axi4_0_awready; 
  assign axi4buf_auto_out_wready = mmio_axi4_0_wready; 
  assign axi4buf_auto_out_bvalid = mmio_axi4_0_bvalid; 
  assign axi4buf_auto_out_bresp = mmio_axi4_0_bresp; 
  assign axi4buf_auto_out_arready = mmio_axi4_0_arready; 
  assign axi4buf_auto_out_rvalid = mmio_axi4_0_rvalid; 
  assign axi4buf_auto_out_rdata = mmio_axi4_0_rdata; 
  assign axi4buf_auto_out_rresp = mmio_axi4_0_rresp; 
  assign axi4buf_auto_out_rlast = mmio_axi4_0_rlast; 
  assign axi4yank_1_clock = clock; 
  assign axi4yank_1_reset = reset; 
  assign axi4yank_1_auto_in_awvalid = axi4deint_auto_out_awvalid; 
  assign axi4yank_1_auto_in_awaddr = axi4deint_auto_out_awaddr; 
  assign axi4yank_1_auto_in_awlen = axi4deint_auto_out_awlen; 
  assign axi4yank_1_auto_in_awsize = axi4deint_auto_out_awsize; 
  assign axi4yank_1_auto_in_awburst = axi4deint_auto_out_awburst; 
  assign axi4yank_1_auto_in_awlock = axi4deint_auto_out_awlock; 
  assign axi4yank_1_auto_in_awcache = axi4deint_auto_out_awcache; 
  assign axi4yank_1_auto_in_awprot = axi4deint_auto_out_awprot; 
  assign axi4yank_1_auto_in_awqos = axi4deint_auto_out_awqos; 
  assign axi4yank_1_auto_in_awuser = axi4deint_auto_out_awuser; 
  assign axi4yank_1_auto_in_awinstret = axi4deint_auto_out_awinstret; 
  assign axi4yank_1_auto_in_wvalid = axi4deint_auto_out_wvalid; 
  assign axi4yank_1_auto_in_wdata = axi4deint_auto_out_wdata; 
  assign axi4yank_1_auto_in_wstrb = axi4deint_auto_out_wstrb; 
  assign axi4yank_1_auto_in_wlast = axi4deint_auto_out_wlast; 
  assign axi4yank_1_auto_in_bready = axi4deint_auto_out_bready; 
  assign axi4yank_1_auto_in_arvalid = axi4deint_auto_out_arvalid; 
  assign axi4yank_1_auto_in_araddr = axi4deint_auto_out_araddr; 
  assign axi4yank_1_auto_in_arlen = axi4deint_auto_out_arlen; 
  assign axi4yank_1_auto_in_arsize = axi4deint_auto_out_arsize; 
  assign axi4yank_1_auto_in_arburst = axi4deint_auto_out_arburst; 
  assign axi4yank_1_auto_in_arlock = axi4deint_auto_out_arlock; 
  assign axi4yank_1_auto_in_arcache = axi4deint_auto_out_arcache; 
  assign axi4yank_1_auto_in_arprot = axi4deint_auto_out_arprot; 
  assign axi4yank_1_auto_in_arqos = axi4deint_auto_out_arqos; 
  assign axi4yank_1_auto_in_aruser = axi4deint_auto_out_aruser; 
  assign axi4yank_1_auto_in_arinstret = axi4deint_auto_out_arinstret; 
  assign axi4yank_1_auto_in_rready = axi4deint_auto_out_rready; 
  assign axi4yank_1_auto_out_awready = axi4buf_auto_in_awready; 
  assign axi4yank_1_auto_out_wready = axi4buf_auto_in_wready; 
  assign axi4yank_1_auto_out_bvalid = axi4buf_auto_in_bvalid; 
  assign axi4yank_1_auto_out_bresp = axi4buf_auto_in_bresp; 
  assign axi4yank_1_auto_out_arready = axi4buf_auto_in_arready; 
  assign axi4yank_1_auto_out_rvalid = axi4buf_auto_in_rvalid; 
  assign axi4yank_1_auto_out_rdata = axi4buf_auto_in_rdata; 
  assign axi4yank_1_auto_out_rresp = axi4buf_auto_in_rresp; 
  assign axi4yank_1_auto_out_rlast = axi4buf_auto_in_rlast; 
  assign axi4deint_clock = clock; 
  assign axi4deint_reset = reset; 
  assign axi4deint_auto_in_awvalid = axi4index_1_auto_out_awvalid; 
  assign axi4deint_auto_in_awaddr = axi4index_1_auto_out_awaddr; 
  assign axi4deint_auto_in_awlen = axi4index_1_auto_out_awlen; 
  assign axi4deint_auto_in_awsize = axi4index_1_auto_out_awsize; 
  assign axi4deint_auto_in_awburst = axi4index_1_auto_out_awburst; 
  assign axi4deint_auto_in_awlock = axi4index_1_auto_out_awlock; 
  assign axi4deint_auto_in_awcache = axi4index_1_auto_out_awcache; 
  assign axi4deint_auto_in_awprot = axi4index_1_auto_out_awprot; 
  assign axi4deint_auto_in_awqos = axi4index_1_auto_out_awqos; 
  assign axi4deint_auto_in_awuser = axi4index_1_auto_out_awuser; 
  assign axi4deint_auto_in_awinstret = axi4index_1_auto_out_awinstret; 
  assign axi4deint_auto_in_wvalid = axi4index_1_auto_out_wvalid; 
  assign axi4deint_auto_in_wdata = axi4index_1_auto_out_wdata; 
  assign axi4deint_auto_in_wstrb = axi4index_1_auto_out_wstrb; 
  assign axi4deint_auto_in_wlast = axi4index_1_auto_out_wlast; 
  assign axi4deint_auto_in_bready = axi4index_1_auto_out_bready; 
  assign axi4deint_auto_in_arvalid = axi4index_1_auto_out_arvalid; 
  assign axi4deint_auto_in_araddr = axi4index_1_auto_out_araddr; 
  assign axi4deint_auto_in_arlen = axi4index_1_auto_out_arlen; 
  assign axi4deint_auto_in_arsize = axi4index_1_auto_out_arsize; 
  assign axi4deint_auto_in_arburst = axi4index_1_auto_out_arburst; 
  assign axi4deint_auto_in_arlock = axi4index_1_auto_out_arlock; 
  assign axi4deint_auto_in_arcache = axi4index_1_auto_out_arcache; 
  assign axi4deint_auto_in_arprot = axi4index_1_auto_out_arprot; 
  assign axi4deint_auto_in_arqos = axi4index_1_auto_out_arqos; 
  assign axi4deint_auto_in_aruser = axi4index_1_auto_out_aruser; 
  assign axi4deint_auto_in_arinstret = axi4index_1_auto_out_arinstret; 
  assign axi4deint_auto_in_rready = axi4index_1_auto_out_rready; 
  assign axi4deint_auto_out_awready = axi4yank_1_auto_in_awready; 
  assign axi4deint_auto_out_wready = axi4yank_1_auto_in_wready; 
  assign axi4deint_auto_out_bvalid = axi4yank_1_auto_in_bvalid; 
  assign axi4deint_auto_out_bresp = axi4yank_1_auto_in_bresp; 
  assign axi4deint_auto_out_buser = axi4yank_1_auto_in_buser; 
  assign axi4deint_auto_out_arready = axi4yank_1_auto_in_arready; 
  assign axi4deint_auto_out_rvalid = axi4yank_1_auto_in_rvalid; 
  assign axi4deint_auto_out_rdata = axi4yank_1_auto_in_rdata; 
  assign axi4deint_auto_out_rresp = axi4yank_1_auto_in_rresp; 
  assign axi4deint_auto_out_ruser = axi4yank_1_auto_in_ruser; 
  assign axi4deint_auto_out_rlast = axi4yank_1_auto_in_rlast; 
  assign axi4index_1_auto_in_awvalid = tl2axi4_1_auto_out_awvalid; 
  assign axi4index_1_auto_in_awid = tl2axi4_1_auto_out_awid; 
  assign axi4index_1_auto_in_awaddr = tl2axi4_1_auto_out_awaddr; 
  assign axi4index_1_auto_in_awlen = tl2axi4_1_auto_out_awlen; 
  assign axi4index_1_auto_in_awsize = tl2axi4_1_auto_out_awsize; 
  assign axi4index_1_auto_in_awburst = tl2axi4_1_auto_out_awburst; 
  assign axi4index_1_auto_in_awlock = tl2axi4_1_auto_out_awlock; 
  assign axi4index_1_auto_in_awcache = tl2axi4_1_auto_out_awcache; 
  assign axi4index_1_auto_in_awprot = tl2axi4_1_auto_out_awprot; 
  assign axi4index_1_auto_in_awqos = tl2axi4_1_auto_out_awqos; 
  assign axi4index_1_auto_in_awuser = tl2axi4_1_auto_out_awuser; 
  assign axi4index_1_auto_in_awinstret = tl2axi4_1_auto_out_awinstret; 
  assign axi4index_1_auto_in_wvalid = tl2axi4_1_auto_out_wvalid; 
  assign axi4index_1_auto_in_wdata = tl2axi4_1_auto_out_wdata; 
  assign axi4index_1_auto_in_wstrb = tl2axi4_1_auto_out_wstrb; 
  assign axi4index_1_auto_in_wlast = tl2axi4_1_auto_out_wlast; 
  assign axi4index_1_auto_in_bready = tl2axi4_1_auto_out_bready; 
  assign axi4index_1_auto_in_arvalid = tl2axi4_1_auto_out_arvalid; 
  assign axi4index_1_auto_in_arid = tl2axi4_1_auto_out_arid; 
  assign axi4index_1_auto_in_araddr = tl2axi4_1_auto_out_araddr; 
  assign axi4index_1_auto_in_arlen = tl2axi4_1_auto_out_arlen; 
  assign axi4index_1_auto_in_arsize = tl2axi4_1_auto_out_arsize; 
  assign axi4index_1_auto_in_arburst = tl2axi4_1_auto_out_arburst; 
  assign axi4index_1_auto_in_arlock = tl2axi4_1_auto_out_arlock; 
  assign axi4index_1_auto_in_arcache = tl2axi4_1_auto_out_arcache; 
  assign axi4index_1_auto_in_arprot = tl2axi4_1_auto_out_arprot; 
  assign axi4index_1_auto_in_arqos = tl2axi4_1_auto_out_arqos; 
  assign axi4index_1_auto_in_aruser = tl2axi4_1_auto_out_aruser; 
  assign axi4index_1_auto_in_arinstret = tl2axi4_1_auto_out_arinstret; 
  assign axi4index_1_auto_in_rready = tl2axi4_1_auto_out_rready; 
  assign axi4index_1_auto_out_awready = axi4deint_auto_in_awready; 
  assign axi4index_1_auto_out_wready = axi4deint_auto_in_wready; 
  assign axi4index_1_auto_out_bvalid = axi4deint_auto_in_bvalid; 
  assign axi4index_1_auto_out_bresp = axi4deint_auto_in_bresp; 
  assign axi4index_1_auto_out_buser = axi4deint_auto_in_buser; 
  assign axi4index_1_auto_out_arready = axi4deint_auto_in_arready; 
  assign axi4index_1_auto_out_rvalid = axi4deint_auto_in_rvalid; 
  assign axi4index_1_auto_out_rdata = axi4deint_auto_in_rdata; 
  assign axi4index_1_auto_out_rresp = axi4deint_auto_in_rresp; 
  assign axi4index_1_auto_out_ruser = axi4deint_auto_in_ruser; 
  assign axi4index_1_auto_out_rlast = axi4deint_auto_in_rlast; 
  assign tl2axi4_1_clock = clock; 
  assign tl2axi4_1_reset = reset; 
  assign tl2axi4_1_auto_in_a_valid = xbar_auto_out_1_a_valid; 
  assign tl2axi4_1_auto_in_a_bits_opcode = xbar_auto_out_1_a_bits_opcode; 
  assign tl2axi4_1_auto_in_a_bits_param = xbar_auto_out_1_a_bits_param; 
  assign tl2axi4_1_auto_in_a_bits_size = xbar_auto_out_1_a_bits_size; 
  assign tl2axi4_1_auto_in_a_bits_source = xbar_auto_out_1_a_bits_source; 
  assign tl2axi4_1_auto_in_a_bits_address = xbar_auto_out_1_a_bits_address; 
  assign tl2axi4_1_auto_in_a_bits_mask = xbar_auto_out_1_a_bits_mask; 
  assign tl2axi4_1_auto_in_a_bits_data = xbar_auto_out_1_a_bits_data; 
  assign tl2axi4_1_auto_in_a_bits_corrupt = xbar_auto_out_1_a_bits_corrupt; 
  assign tl2axi4_1_auto_in_d_ready = xbar_auto_out_1_d_ready; 
  assign tl2axi4_1_auto_out_awready = axi4index_1_auto_in_awready; 
  assign tl2axi4_1_auto_out_wready = axi4index_1_auto_in_wready; 
  assign tl2axi4_1_auto_out_bvalid = axi4index_1_auto_in_bvalid; 
  assign tl2axi4_1_auto_out_bid = axi4index_1_auto_in_bid; 
  assign tl2axi4_1_auto_out_bresp = axi4index_1_auto_in_bresp; 
  assign tl2axi4_1_auto_out_buser = axi4index_1_auto_in_buser; 
  assign tl2axi4_1_auto_out_arready = axi4index_1_auto_in_arready; 
  assign tl2axi4_1_auto_out_rvalid = axi4index_1_auto_in_rvalid; 
  assign tl2axi4_1_auto_out_rid = axi4index_1_auto_in_rid; 
  assign tl2axi4_1_auto_out_rdata = axi4index_1_auto_in_rdata; 
  assign tl2axi4_1_auto_out_rresp = axi4index_1_auto_in_rresp; 
  assign tl2axi4_1_auto_out_ruser = axi4index_1_auto_in_ruser; 
  assign tl2axi4_1_auto_out_rlast = axi4index_1_auto_in_rlast; 
  assign fixer_clock = clock; 
  assign fixer_reset = reset; 
  assign fixer_auto_in_a_valid = widget_auto_out_a_valid; 
  assign fixer_auto_in_a_bits_opcode = widget_auto_out_a_bits_opcode; 
  assign fixer_auto_in_a_bits_param = widget_auto_out_a_bits_param; 
  assign fixer_auto_in_a_bits_size = widget_auto_out_a_bits_size; 
  assign fixer_auto_in_a_bits_source = widget_auto_out_a_bits_source; 
  assign fixer_auto_in_a_bits_address = widget_auto_out_a_bits_address; 
  assign fixer_auto_in_a_bits_mask = widget_auto_out_a_bits_mask; 
  assign fixer_auto_in_a_bits_data = widget_auto_out_a_bits_data; 
  assign fixer_auto_in_a_bits_corrupt = widget_auto_out_a_bits_corrupt; 
  assign fixer_auto_in_d_ready = widget_auto_out_d_ready; 
  assign fixer_auto_out_a_ready = xbar_1_auto_in_a_ready; 
  assign fixer_auto_out_d_valid = xbar_1_auto_in_d_valid; 
  assign fixer_auto_out_d_bits_opcode = xbar_1_auto_in_d_bits_opcode; 
  assign fixer_auto_out_d_bits_param = xbar_1_auto_in_d_bits_param; 
  assign fixer_auto_out_d_bits_size = xbar_1_auto_in_d_bits_size; 
  assign fixer_auto_out_d_bits_source = xbar_1_auto_in_d_bits_source; 
  assign fixer_auto_out_d_bits_sink = xbar_1_auto_in_d_bits_sink; 
  assign fixer_auto_out_d_bits_denied = xbar_1_auto_in_d_bits_denied; 
  assign fixer_auto_out_d_bits_data = xbar_1_auto_in_d_bits_data; 
  assign fixer_auto_out_d_bits_corrupt = xbar_1_auto_in_d_bits_corrupt; 
  assign widget_clock = clock; 
  assign widget_reset = reset; 
  assign widget_auto_in_a_valid = axi42tl_auto_out_a_valid; 
  assign widget_auto_in_a_bits_opcode = axi42tl_auto_out_a_bits_opcode; 
  assign widget_auto_in_a_bits_param = axi42tl_auto_out_a_bits_param; 
  assign widget_auto_in_a_bits_size = axi42tl_auto_out_a_bits_size; 
  assign widget_auto_in_a_bits_source = axi42tl_auto_out_a_bits_source; 
  assign widget_auto_in_a_bits_address = axi42tl_auto_out_a_bits_address; 
  assign widget_auto_in_a_bits_mask = axi42tl_auto_out_a_bits_mask; 
  assign widget_auto_in_a_bits_data = axi42tl_auto_out_a_bits_data; 
  assign widget_auto_in_a_bits_corrupt = axi42tl_auto_out_a_bits_corrupt; 
  assign widget_auto_in_d_ready = axi42tl_auto_out_d_ready; 
  assign widget_auto_out_a_ready = fixer_auto_in_a_ready; 
  assign widget_auto_out_d_valid = fixer_auto_in_d_valid; 
  assign widget_auto_out_d_bits_opcode = fixer_auto_in_d_bits_opcode; 
  assign widget_auto_out_d_bits_param = fixer_auto_in_d_bits_param; 
  assign widget_auto_out_d_bits_size = fixer_auto_in_d_bits_size; 
  assign widget_auto_out_d_bits_source = fixer_auto_in_d_bits_source; 
  assign widget_auto_out_d_bits_sink = fixer_auto_in_d_bits_sink; 
  assign widget_auto_out_d_bits_denied = fixer_auto_in_d_bits_denied; 
  assign widget_auto_out_d_bits_data = fixer_auto_in_d_bits_data; 
  assign widget_auto_out_d_bits_corrupt = fixer_auto_in_d_bits_corrupt; 
  assign axi42tl_clock = clock; 
  assign axi42tl_reset = reset; 
  assign axi42tl_auto_in_awvalid = axi4yank_2_auto_out_awvalid; 
  assign axi42tl_auto_in_awid = axi4yank_2_auto_out_awid; 
  assign axi42tl_auto_in_awaddr = axi4yank_2_auto_out_awaddr; 
  assign axi42tl_auto_in_awlen = axi4yank_2_auto_out_awlen; 
  assign axi42tl_auto_in_awsize = axi4yank_2_auto_out_awsize; 
  assign axi42tl_auto_in_wvalid = axi4yank_2_auto_out_wvalid; 
  assign axi42tl_auto_in_wdata = axi4yank_2_auto_out_wdata; 
  assign axi42tl_auto_in_wstrb = axi4yank_2_auto_out_wstrb; 
  assign axi42tl_auto_in_wlast = axi4yank_2_auto_out_wlast; 
  assign axi42tl_auto_in_bready = axi4yank_2_auto_out_bready; 
  assign axi42tl_auto_in_arvalid = axi4yank_2_auto_out_arvalid; 
  assign axi42tl_auto_in_arid = axi4yank_2_auto_out_arid; 
  assign axi42tl_auto_in_araddr = axi4yank_2_auto_out_araddr; 
  assign axi42tl_auto_in_arlen = axi4yank_2_auto_out_arlen; 
  assign axi42tl_auto_in_arsize = axi4yank_2_auto_out_arsize; 
  assign axi42tl_auto_in_rready = axi4yank_2_auto_out_rready; 
  assign axi42tl_auto_out_a_ready = widget_auto_in_a_ready; 
  assign axi42tl_auto_out_d_valid = widget_auto_in_d_valid; 
  assign axi42tl_auto_out_d_bits_opcode = widget_auto_in_d_bits_opcode; 
  assign axi42tl_auto_out_d_bits_size = widget_auto_in_d_bits_size; 
  assign axi42tl_auto_out_d_bits_source = widget_auto_in_d_bits_source; 
  assign axi42tl_auto_out_d_bits_denied = widget_auto_in_d_bits_denied; 
  assign axi42tl_auto_out_d_bits_data = widget_auto_in_d_bits_data; 
  assign axi42tl_auto_out_d_bits_corrupt = widget_auto_in_d_bits_corrupt; 
  assign axi4yank_2_clock = clock; 
  assign axi4yank_2_reset = reset; 
  assign axi4yank_2_auto_in_awvalid = axi4frag_auto_out_awvalid; 
  assign axi4yank_2_auto_in_awid = axi4frag_auto_out_awid; 
  assign axi4yank_2_auto_in_awaddr = axi4frag_auto_out_awaddr; 
  assign axi4yank_2_auto_in_awlen = axi4frag_auto_out_awlen; 
  assign axi4yank_2_auto_in_awsize = axi4frag_auto_out_awsize; 
  assign axi4yank_2_auto_in_awuser = axi4frag_auto_out_awuser; 
  assign axi4yank_2_auto_in_wvalid = axi4frag_auto_out_wvalid; 
  assign axi4yank_2_auto_in_wdata = axi4frag_auto_out_wdata; 
  assign axi4yank_2_auto_in_wstrb = axi4frag_auto_out_wstrb; 
  assign axi4yank_2_auto_in_wlast = axi4frag_auto_out_wlast; 
  assign axi4yank_2_auto_in_bready = axi4frag_auto_out_bready; 
  assign axi4yank_2_auto_in_arvalid = axi4frag_auto_out_arvalid; 
  assign axi4yank_2_auto_in_arid = axi4frag_auto_out_arid; 
  assign axi4yank_2_auto_in_araddr = axi4frag_auto_out_araddr; 
  assign axi4yank_2_auto_in_arlen = axi4frag_auto_out_arlen; 
  assign axi4yank_2_auto_in_arsize = axi4frag_auto_out_arsize; 
  assign axi4yank_2_auto_in_aruser = axi4frag_auto_out_aruser; 
  assign axi4yank_2_auto_in_rready = axi4frag_auto_out_rready; 
  assign axi4yank_2_auto_out_awready = axi42tl_auto_in_awready; 
  assign axi4yank_2_auto_out_wready = axi42tl_auto_in_wready; 
  assign axi4yank_2_auto_out_bvalid = axi42tl_auto_in_bvalid; 
  assign axi4yank_2_auto_out_bid = axi42tl_auto_in_bid; 
  assign axi4yank_2_auto_out_bresp = axi42tl_auto_in_bresp; 
  assign axi4yank_2_auto_out_arready = axi42tl_auto_in_arready; 
  assign axi4yank_2_auto_out_rvalid = axi42tl_auto_in_rvalid; 
  assign axi4yank_2_auto_out_rid = axi42tl_auto_in_rid; 
  assign axi4yank_2_auto_out_rdata = axi42tl_auto_in_rdata; 
  assign axi4yank_2_auto_out_rresp = axi42tl_auto_in_rresp; 
  assign axi4yank_2_auto_out_rlast = axi42tl_auto_in_rlast; 
  assign axi4frag_clock = clock; 
  assign axi4frag_reset = reset; 
  assign axi4frag_auto_in_awvalid = axi4index_2_auto_out_awvalid; 
  assign axi4frag_auto_in_awid = axi4index_2_auto_out_awid; 
  assign axi4frag_auto_in_awaddr = axi4index_2_auto_out_awaddr; 
  assign axi4frag_auto_in_awlen = axi4index_2_auto_out_awlen; 
  assign axi4frag_auto_in_awsize = axi4index_2_auto_out_awsize; 
  assign axi4frag_auto_in_awburst = axi4index_2_auto_out_awburst; 
  assign axi4frag_auto_in_awuser = axi4index_2_auto_out_awuser; 
  assign axi4frag_auto_in_wvalid = axi4index_2_auto_out_wvalid; 
  assign axi4frag_auto_in_wdata = axi4index_2_auto_out_wdata; 
  assign axi4frag_auto_in_wstrb = axi4index_2_auto_out_wstrb; 
  assign axi4frag_auto_in_wlast = axi4index_2_auto_out_wlast; 
  assign axi4frag_auto_in_bready = axi4index_2_auto_out_bready; 
  assign axi4frag_auto_in_arvalid = axi4index_2_auto_out_arvalid; 
  assign axi4frag_auto_in_arid = axi4index_2_auto_out_arid; 
  assign axi4frag_auto_in_araddr = axi4index_2_auto_out_araddr; 
  assign axi4frag_auto_in_arlen = axi4index_2_auto_out_arlen; 
  assign axi4frag_auto_in_arsize = axi4index_2_auto_out_arsize; 
  assign axi4frag_auto_in_arburst = axi4index_2_auto_out_arburst; 
  assign axi4frag_auto_in_aruser = axi4index_2_auto_out_aruser; 
  assign axi4frag_auto_in_rready = axi4index_2_auto_out_rready; 
  assign axi4frag_auto_out_awready = axi4yank_2_auto_in_awready; 
  assign axi4frag_auto_out_wready = axi4yank_2_auto_in_wready; 
  assign axi4frag_auto_out_bvalid = axi4yank_2_auto_in_bvalid; 
  assign axi4frag_auto_out_bid = axi4yank_2_auto_in_bid; 
  assign axi4frag_auto_out_bresp = axi4yank_2_auto_in_bresp; 
  assign axi4frag_auto_out_buser = axi4yank_2_auto_in_buser; 
  assign axi4frag_auto_out_arready = axi4yank_2_auto_in_arready; 
  assign axi4frag_auto_out_rvalid = axi4yank_2_auto_in_rvalid; 
  assign axi4frag_auto_out_rid = axi4yank_2_auto_in_rid; 
  assign axi4frag_auto_out_rdata = axi4yank_2_auto_in_rdata; 
  assign axi4frag_auto_out_rresp = axi4yank_2_auto_in_rresp; 
  assign axi4frag_auto_out_ruser = axi4yank_2_auto_in_ruser; 
  assign axi4frag_auto_out_rlast = axi4yank_2_auto_in_rlast; 
  assign axi4index_2_auto_in_awvalid = l2_frontend_bus_axi4_0_awvalid; 
  assign axi4index_2_auto_in_awid = l2_frontend_bus_axi4_0_awid; 
  assign axi4index_2_auto_in_awaddr = l2_frontend_bus_axi4_0_awaddr; 
  assign axi4index_2_auto_in_awlen = l2_frontend_bus_axi4_0_awlen; 
  assign axi4index_2_auto_in_awsize = l2_frontend_bus_axi4_0_awsize; 
  assign axi4index_2_auto_in_awburst = l2_frontend_bus_axi4_0_awburst; 
  assign axi4index_2_auto_in_wvalid = l2_frontend_bus_axi4_0_wvalid; 
  assign axi4index_2_auto_in_wdata = l2_frontend_bus_axi4_0_wdata; 
  assign axi4index_2_auto_in_wstrb = l2_frontend_bus_axi4_0_wstrb; 
  assign axi4index_2_auto_in_wlast = l2_frontend_bus_axi4_0_wlast; 
  assign axi4index_2_auto_in_bready = l2_frontend_bus_axi4_0_bready; 
  assign axi4index_2_auto_in_arvalid = l2_frontend_bus_axi4_0_arvalid; 
  assign axi4index_2_auto_in_arid = l2_frontend_bus_axi4_0_arid; 
  assign axi4index_2_auto_in_araddr = l2_frontend_bus_axi4_0_araddr; 
  assign axi4index_2_auto_in_arlen = l2_frontend_bus_axi4_0_arlen; 
  assign axi4index_2_auto_in_arsize = l2_frontend_bus_axi4_0_arsize; 
  assign axi4index_2_auto_in_arburst = l2_frontend_bus_axi4_0_arburst; 
  assign axi4index_2_auto_in_rready = l2_frontend_bus_axi4_0_rready; 
  assign axi4index_2_auto_out_awready = axi4frag_auto_in_awready; 
  assign axi4index_2_auto_out_wready = axi4frag_auto_in_wready; 
  assign axi4index_2_auto_out_bvalid = axi4frag_auto_in_bvalid; 
  assign axi4index_2_auto_out_bid = axi4frag_auto_in_bid; 
  assign axi4index_2_auto_out_bresp = axi4frag_auto_in_bresp; 
  assign axi4index_2_auto_out_buser = axi4frag_auto_in_buser; 
  assign axi4index_2_auto_out_arready = axi4frag_auto_in_arready; 
  assign axi4index_2_auto_out_rvalid = axi4frag_auto_in_rvalid; 
  assign axi4index_2_auto_out_rid = axi4frag_auto_in_rid; 
  assign axi4index_2_auto_out_rdata = axi4frag_auto_in_rdata; 
  assign axi4index_2_auto_out_rresp = axi4frag_auto_in_rresp; 
  assign axi4index_2_auto_out_ruser = axi4frag_auto_in_ruser; 
  assign axi4index_2_auto_out_rlast = axi4frag_auto_in_rlast; 
  assign err_clock = clock; 
  assign err_reset = reset; 
  assign err_auto_in_a_valid = widget_2_auto_out_a_valid; 
  assign err_auto_in_a_bits_opcode = widget_2_auto_out_a_bits_opcode; 
  assign err_auto_in_a_bits_param = widget_2_auto_out_a_bits_param; 
  assign err_auto_in_a_bits_size = widget_2_auto_out_a_bits_size; 
  assign err_auto_in_a_bits_source = widget_2_auto_out_a_bits_source; 
  assign err_auto_in_a_bits_address = widget_2_auto_out_a_bits_address; 
  assign err_auto_in_a_bits_mask = widget_2_auto_out_a_bits_mask; 
  assign err_auto_in_a_bits_corrupt = widget_2_auto_out_a_bits_corrupt; 
  assign err_auto_in_c_valid = widget_2_auto_out_c_valid; 
  assign err_auto_in_c_bits_opcode = widget_2_auto_out_c_bits_opcode; 
  assign err_auto_in_c_bits_param = widget_2_auto_out_c_bits_param; 
  assign err_auto_in_c_bits_size = widget_2_auto_out_c_bits_size; 
  assign err_auto_in_c_bits_source = widget_2_auto_out_c_bits_source; 
  assign err_auto_in_c_bits_address = widget_2_auto_out_c_bits_address; 
  assign err_auto_in_c_bits_corrupt = widget_2_auto_out_c_bits_corrupt; 
  assign err_auto_in_d_ready = widget_2_auto_out_d_ready; 
  assign err_auto_in_e_valid = widget_2_auto_out_e_valid; 
  assign atomics_clock = clock; 
  assign atomics_reset = reset; 
  assign atomics_auto_in_a_valid = fixer_1_auto_out_a_valid; 
  assign atomics_auto_in_a_bits_opcode = fixer_1_auto_out_a_bits_opcode; 
  assign atomics_auto_in_a_bits_param = fixer_1_auto_out_a_bits_param; 
  assign atomics_auto_in_a_bits_size = fixer_1_auto_out_a_bits_size; 
  assign atomics_auto_in_a_bits_source = fixer_1_auto_out_a_bits_source; 
  assign atomics_auto_in_a_bits_address = fixer_1_auto_out_a_bits_address; 
  assign atomics_auto_in_a_bits_mask = fixer_1_auto_out_a_bits_mask; 
  assign atomics_auto_in_a_bits_data = fixer_1_auto_out_a_bits_data; 
  assign atomics_auto_in_c_valid = fixer_1_auto_out_c_valid; 
  assign atomics_auto_in_c_bits_opcode = fixer_1_auto_out_c_bits_opcode; 
  assign atomics_auto_in_c_bits_param = fixer_1_auto_out_c_bits_param; 
  assign atomics_auto_in_c_bits_size = fixer_1_auto_out_c_bits_size; 
  assign atomics_auto_in_c_bits_source = fixer_1_auto_out_c_bits_source; 
  assign atomics_auto_in_c_bits_address = fixer_1_auto_out_c_bits_address; 
  assign atomics_auto_in_c_bits_corrupt = fixer_1_auto_out_c_bits_corrupt; 
  assign atomics_auto_in_d_ready = fixer_1_auto_out_d_ready; 
  assign atomics_auto_in_e_valid = fixer_1_auto_out_e_valid; 
  assign atomics_auto_in_e_bits_sink = fixer_1_auto_out_e_bits_sink; 
  assign atomics_auto_out_a_ready = xbar_auto_in_a_ready; 
  assign atomics_auto_out_c_ready = xbar_auto_in_c_ready; 
  assign atomics_auto_out_d_valid = xbar_auto_in_d_valid; 
  assign atomics_auto_out_d_bits_opcode = xbar_auto_in_d_bits_opcode; 
  assign atomics_auto_out_d_bits_param = xbar_auto_in_d_bits_param; 
  assign atomics_auto_out_d_bits_size = xbar_auto_in_d_bits_size; 
  assign atomics_auto_out_d_bits_source = xbar_auto_in_d_bits_source; 
  assign atomics_auto_out_d_bits_sink = xbar_auto_in_d_bits_sink; 
  assign atomics_auto_out_d_bits_denied = xbar_auto_in_d_bits_denied; 
  assign atomics_auto_out_d_bits_data = xbar_auto_in_d_bits_data; 
  assign atomics_auto_out_d_bits_corrupt = xbar_auto_in_d_bits_corrupt; 
  assign atomics_auto_out_e_ready = xbar_auto_in_e_ready; 
  assign fixer_1_clock = clock; 
  assign fixer_1_reset = reset; 
  assign fixer_1_auto_in_a_valid = hints_auto_out_a_valid; 
  assign fixer_1_auto_in_a_bits_opcode = hints_auto_out_a_bits_opcode; 
  assign fixer_1_auto_in_a_bits_param = hints_auto_out_a_bits_param; 
  assign fixer_1_auto_in_a_bits_size = hints_auto_out_a_bits_size; 
  assign fixer_1_auto_in_a_bits_source = hints_auto_out_a_bits_source; 
  assign fixer_1_auto_in_a_bits_address = hints_auto_out_a_bits_address; 
  assign fixer_1_auto_in_a_bits_mask = hints_auto_out_a_bits_mask; 
  assign fixer_1_auto_in_a_bits_data = hints_auto_out_a_bits_data; 
  assign fixer_1_auto_in_c_valid = hints_auto_out_c_valid; 
  assign fixer_1_auto_in_c_bits_opcode = hints_auto_out_c_bits_opcode; 
  assign fixer_1_auto_in_c_bits_param = hints_auto_out_c_bits_param; 
  assign fixer_1_auto_in_c_bits_size = hints_auto_out_c_bits_size; 
  assign fixer_1_auto_in_c_bits_source = hints_auto_out_c_bits_source; 
  assign fixer_1_auto_in_c_bits_address = hints_auto_out_c_bits_address; 
  assign fixer_1_auto_in_c_bits_corrupt = hints_auto_out_c_bits_corrupt; 
  assign fixer_1_auto_in_d_ready = hints_auto_out_d_ready; 
  assign fixer_1_auto_in_e_valid = hints_auto_out_e_valid; 
  assign fixer_1_auto_in_e_bits_sink = hints_auto_out_e_bits_sink; 
  assign fixer_1_auto_out_a_ready = atomics_auto_in_a_ready; 
  assign fixer_1_auto_out_c_ready = atomics_auto_in_c_ready; 
  assign fixer_1_auto_out_d_valid = atomics_auto_in_d_valid; 
  assign fixer_1_auto_out_d_bits_opcode = atomics_auto_in_d_bits_opcode; 
  assign fixer_1_auto_out_d_bits_param = atomics_auto_in_d_bits_param; 
  assign fixer_1_auto_out_d_bits_size = atomics_auto_in_d_bits_size; 
  assign fixer_1_auto_out_d_bits_source = atomics_auto_in_d_bits_source; 
  assign fixer_1_auto_out_d_bits_sink = atomics_auto_in_d_bits_sink; 
  assign fixer_1_auto_out_d_bits_denied = atomics_auto_in_d_bits_denied; 
  assign fixer_1_auto_out_d_bits_data = atomics_auto_in_d_bits_data; 
  assign fixer_1_auto_out_d_bits_corrupt = atomics_auto_in_d_bits_corrupt; 
  assign fixer_1_auto_out_e_ready = atomics_auto_in_e_ready; 
  assign hints_clock = clock; 
  assign hints_reset = reset; 
  assign hints_auto_in_a_valid = widget_1_auto_out_a_valid; 
  assign hints_auto_in_a_bits_opcode = widget_1_auto_out_a_bits_opcode; 
  assign hints_auto_in_a_bits_param = widget_1_auto_out_a_bits_param; 
  assign hints_auto_in_a_bits_size = widget_1_auto_out_a_bits_size; 
  assign hints_auto_in_a_bits_source = widget_1_auto_out_a_bits_source; 
  assign hints_auto_in_a_bits_address = widget_1_auto_out_a_bits_address; 
  assign hints_auto_in_a_bits_mask = widget_1_auto_out_a_bits_mask; 
  assign hints_auto_in_a_bits_data = widget_1_auto_out_a_bits_data; 
  assign hints_auto_in_c_valid = widget_1_auto_out_c_valid; 
  assign hints_auto_in_c_bits_opcode = widget_1_auto_out_c_bits_opcode; 
  assign hints_auto_in_c_bits_param = widget_1_auto_out_c_bits_param; 
  assign hints_auto_in_c_bits_size = widget_1_auto_out_c_bits_size; 
  assign hints_auto_in_c_bits_source = widget_1_auto_out_c_bits_source; 
  assign hints_auto_in_c_bits_address = widget_1_auto_out_c_bits_address; 
  assign hints_auto_in_c_bits_corrupt = widget_1_auto_out_c_bits_corrupt; 
  assign hints_auto_in_d_ready = widget_1_auto_out_d_ready; 
  assign hints_auto_in_e_valid = widget_1_auto_out_e_valid; 
  assign hints_auto_in_e_bits_sink = widget_1_auto_out_e_bits_sink; 
  assign hints_auto_out_a_ready = fixer_1_auto_in_a_ready; 
  assign hints_auto_out_c_ready = fixer_1_auto_in_c_ready; 
  assign hints_auto_out_d_valid = fixer_1_auto_in_d_valid; 
  assign hints_auto_out_d_bits_opcode = fixer_1_auto_in_d_bits_opcode; 
  assign hints_auto_out_d_bits_param = fixer_1_auto_in_d_bits_param; 
  assign hints_auto_out_d_bits_size = fixer_1_auto_in_d_bits_size; 
  assign hints_auto_out_d_bits_source = fixer_1_auto_in_d_bits_source; 
  assign hints_auto_out_d_bits_sink = fixer_1_auto_in_d_bits_sink; 
  assign hints_auto_out_d_bits_denied = fixer_1_auto_in_d_bits_denied; 
  assign hints_auto_out_d_bits_data = fixer_1_auto_in_d_bits_data; 
  assign hints_auto_out_d_bits_corrupt = fixer_1_auto_in_d_bits_corrupt; 
  assign hints_auto_out_e_ready = fixer_1_auto_in_e_ready; 
  assign widget_1_clock = clock; 
  assign widget_1_reset = reset; 
  assign widget_1_auto_in_a_valid = chiplink_auto_mbypass_out_a_valid; 
  assign widget_1_auto_in_a_bits_opcode = chiplink_auto_mbypass_out_a_bits_opcode; 
  assign widget_1_auto_in_a_bits_param = chiplink_auto_mbypass_out_a_bits_param; 
  assign widget_1_auto_in_a_bits_size = chiplink_auto_mbypass_out_a_bits_size; 
  assign widget_1_auto_in_a_bits_source = chiplink_auto_mbypass_out_a_bits_source; 
  assign widget_1_auto_in_a_bits_address = chiplink_auto_mbypass_out_a_bits_address; 
  assign widget_1_auto_in_a_bits_mask = chiplink_auto_mbypass_out_a_bits_mask; 
  assign widget_1_auto_in_a_bits_data = chiplink_auto_mbypass_out_a_bits_data; 
  assign widget_1_auto_in_c_valid = chiplink_auto_mbypass_out_c_valid; 
  assign widget_1_auto_in_c_bits_opcode = chiplink_auto_mbypass_out_c_bits_opcode; 
  assign widget_1_auto_in_c_bits_param = chiplink_auto_mbypass_out_c_bits_param; 
  assign widget_1_auto_in_c_bits_size = chiplink_auto_mbypass_out_c_bits_size; 
  assign widget_1_auto_in_c_bits_source = chiplink_auto_mbypass_out_c_bits_source; 
  assign widget_1_auto_in_c_bits_address = chiplink_auto_mbypass_out_c_bits_address; 
  assign widget_1_auto_in_c_bits_corrupt = chiplink_auto_mbypass_out_c_bits_corrupt; 
  assign widget_1_auto_in_d_ready = chiplink_auto_mbypass_out_d_ready; 
  assign widget_1_auto_in_e_valid = chiplink_auto_mbypass_out_e_valid; 
  assign widget_1_auto_in_e_bits_sink = chiplink_auto_mbypass_out_e_bits_sink; 
  assign widget_1_auto_out_a_ready = hints_auto_in_a_ready; 
  assign widget_1_auto_out_c_ready = hints_auto_in_c_ready; 
  assign widget_1_auto_out_d_valid = hints_auto_in_d_valid; 
  assign widget_1_auto_out_d_bits_opcode = hints_auto_in_d_bits_opcode; 
  assign widget_1_auto_out_d_bits_param = hints_auto_in_d_bits_param; 
  assign widget_1_auto_out_d_bits_size = hints_auto_in_d_bits_size; 
  assign widget_1_auto_out_d_bits_source = hints_auto_in_d_bits_source; 
  assign widget_1_auto_out_d_bits_sink = hints_auto_in_d_bits_sink; 
  assign widget_1_auto_out_d_bits_denied = hints_auto_in_d_bits_denied; 
  assign widget_1_auto_out_d_bits_data = hints_auto_in_d_bits_data; 
  assign widget_1_auto_out_d_bits_corrupt = hints_auto_in_d_bits_corrupt; 
  assign widget_1_auto_out_e_ready = hints_auto_in_e_ready; 
  assign widget_2_clock = clock; 
  assign widget_2_reset = reset; 
  assign widget_2_auto_in_a_valid = xbar_auto_out_2_a_valid; 
  assign widget_2_auto_in_a_bits_opcode = xbar_auto_out_2_a_bits_opcode; 
  assign widget_2_auto_in_a_bits_param = xbar_auto_out_2_a_bits_param; 
  assign widget_2_auto_in_a_bits_size = xbar_auto_out_2_a_bits_size; 
  assign widget_2_auto_in_a_bits_source = xbar_auto_out_2_a_bits_source; 
  assign widget_2_auto_in_a_bits_address = xbar_auto_out_2_a_bits_address; 
  assign widget_2_auto_in_a_bits_mask = xbar_auto_out_2_a_bits_mask; 
  assign widget_2_auto_in_a_bits_corrupt = xbar_auto_out_2_a_bits_corrupt; 
  assign widget_2_auto_in_c_valid = xbar_auto_out_2_c_valid; 
  assign widget_2_auto_in_c_bits_opcode = xbar_auto_out_2_c_bits_opcode; 
  assign widget_2_auto_in_c_bits_param = xbar_auto_out_2_c_bits_param; 
  assign widget_2_auto_in_c_bits_size = xbar_auto_out_2_c_bits_size; 
  assign widget_2_auto_in_c_bits_source = xbar_auto_out_2_c_bits_source; 
  assign widget_2_auto_in_c_bits_address = xbar_auto_out_2_c_bits_address; 
  assign widget_2_auto_in_c_bits_corrupt = xbar_auto_out_2_c_bits_corrupt; 
  assign widget_2_auto_in_d_ready = xbar_auto_out_2_d_ready; 
  assign widget_2_auto_in_e_valid = xbar_auto_out_2_e_valid; 
  assign widget_2_auto_out_a_ready = err_auto_in_a_ready; 
  assign widget_2_auto_out_c_ready = err_auto_in_c_ready; 
  assign widget_2_auto_out_d_valid = err_auto_in_d_valid; 
  assign widget_2_auto_out_d_bits_opcode = err_auto_in_d_bits_opcode; 
  assign widget_2_auto_out_d_bits_param = err_auto_in_d_bits_param; 
  assign widget_2_auto_out_d_bits_size = err_auto_in_d_bits_size; 
  assign widget_2_auto_out_d_bits_source = err_auto_in_d_bits_source; 
  assign widget_2_auto_out_d_bits_sink = err_auto_in_d_bits_sink; 
  assign widget_2_auto_out_d_bits_denied = err_auto_in_d_bits_denied; 
  assign widget_2_auto_out_d_bits_data = err_auto_in_d_bits_data; 
  assign widget_2_auto_out_d_bits_corrupt = err_auto_in_d_bits_corrupt; 
endmodule
module dual_ChipLink( 
  input         clock, 
  input         reset, 
  input         auto_mbypass_out_a_ready, 
  output        auto_mbypass_out_a_valid, 
  output [2:0]  auto_mbypass_out_a_bits_opcode, 
  output [2:0]  auto_mbypass_out_a_bits_param, 
  output [3:0]  auto_mbypass_out_a_bits_size, 
  output [5:0]  auto_mbypass_out_a_bits_source, 
  output [31:0] auto_mbypass_out_a_bits_address, 
  output [3:0]  auto_mbypass_out_a_bits_mask, 
  output [31:0] auto_mbypass_out_a_bits_data, 
  input         auto_mbypass_out_c_ready, 
  output        auto_mbypass_out_c_valid, 
  output [2:0]  auto_mbypass_out_c_bits_opcode, 
  output [2:0]  auto_mbypass_out_c_bits_param, 
  output [3:0]  auto_mbypass_out_c_bits_size, 
  output [5:0]  auto_mbypass_out_c_bits_source, 
  output [31:0] auto_mbypass_out_c_bits_address, 
  output        auto_mbypass_out_c_bits_corrupt, 
  output        auto_mbypass_out_d_ready, 
  input         auto_mbypass_out_d_valid, 
  input  [2:0]  auto_mbypass_out_d_bits_opcode, 
  input  [1:0]  auto_mbypass_out_d_bits_param, 
  input  [3:0]  auto_mbypass_out_d_bits_size, 
  input  [5:0]  auto_mbypass_out_d_bits_source, 
  input         auto_mbypass_out_d_bits_sink, 
  input         auto_mbypass_out_d_bits_denied, 
  input  [31:0] auto_mbypass_out_d_bits_data, 
  input         auto_mbypass_out_d_bits_corrupt, 
  input         auto_mbypass_out_e_ready, 
  output        auto_mbypass_out_e_valid, 
  output        auto_mbypass_out_e_bits_sink, 
  output        auto_sbypass_node_in_in_a_ready, 
  input         auto_sbypass_node_in_in_a_valid, 
  input  [2:0]  auto_sbypass_node_in_in_a_bits_opcode, 
  input  [2:0]  auto_sbypass_node_in_in_a_bits_param, 
  input  [2:0]  auto_sbypass_node_in_in_a_bits_size, 
  input  [2:0]  auto_sbypass_node_in_in_a_bits_source, 
  input  [31:0] auto_sbypass_node_in_in_a_bits_address, 
  input  [3:0]  auto_sbypass_node_in_in_a_bits_mask, 
  input  [31:0] auto_sbypass_node_in_in_a_bits_data, 
  input         auto_sbypass_node_in_in_a_bits_corrupt, 
  input         auto_sbypass_node_in_in_d_ready, 
  output        auto_sbypass_node_in_in_d_valid, 
  output [2:0]  auto_sbypass_node_in_in_d_bits_opcode, 
  output [1:0]  auto_sbypass_node_in_in_d_bits_param, 
  output [2:0]  auto_sbypass_node_in_in_d_bits_size, 
  output [2:0]  auto_sbypass_node_in_in_d_bits_source, 
  output [4:0]  auto_sbypass_node_in_in_d_bits_sink, 
  output        auto_sbypass_node_in_in_d_bits_denied, 
  output [31:0] auto_sbypass_node_in_in_d_bits_data, 
  output        auto_sbypass_node_in_in_d_bits_corrupt, 
  output        auto_io_out_c2b_clk, 
  output        auto_io_out_c2b_rst, 
  output        auto_io_out_c2b_send, 
  output [31:0] auto_io_out_c2b_data, 
  input         auto_io_out_b2c_clk, 
  input         auto_io_out_b2c_rst, 
  input         auto_io_out_b2c_send, 
  input  [31:0] auto_io_out_b2c_data 
);
  wire  sbypass_clock; 
  wire  sbypass_reset; 
  wire  sbypass_auto_node_out_out_a_ready; 
  wire  sbypass_auto_node_out_out_a_valid; 
  wire [2:0] sbypass_auto_node_out_out_a_bits_opcode; 
  wire [2:0] sbypass_auto_node_out_out_a_bits_param; 
  wire [2:0] sbypass_auto_node_out_out_a_bits_size; 
  wire [2:0] sbypass_auto_node_out_out_a_bits_source; 
  wire [31:0] sbypass_auto_node_out_out_a_bits_address; 
  wire [3:0] sbypass_auto_node_out_out_a_bits_mask; 
  wire [31:0] sbypass_auto_node_out_out_a_bits_data; 
  wire  sbypass_auto_node_out_out_a_bits_corrupt; 
  wire  sbypass_auto_node_out_out_d_ready; 
  wire  sbypass_auto_node_out_out_d_valid; 
  wire [2:0] sbypass_auto_node_out_out_d_bits_opcode; 
  wire [1:0] sbypass_auto_node_out_out_d_bits_param; 
  wire [2:0] sbypass_auto_node_out_out_d_bits_size; 
  wire [2:0] sbypass_auto_node_out_out_d_bits_source; 
  wire [4:0] sbypass_auto_node_out_out_d_bits_sink; 
  wire  sbypass_auto_node_out_out_d_bits_denied; 
  wire [31:0] sbypass_auto_node_out_out_d_bits_data; 
  wire  sbypass_auto_node_out_out_d_bits_corrupt; 
  wire  sbypass_auto_node_in_in_a_ready; 
  wire  sbypass_auto_node_in_in_a_valid; 
  wire [2:0] sbypass_auto_node_in_in_a_bits_opcode; 
  wire [2:0] sbypass_auto_node_in_in_a_bits_param; 
  wire [2:0] sbypass_auto_node_in_in_a_bits_size; 
  wire [2:0] sbypass_auto_node_in_in_a_bits_source; 
  wire [31:0] sbypass_auto_node_in_in_a_bits_address; 
  wire [3:0] sbypass_auto_node_in_in_a_bits_mask; 
  wire [31:0] sbypass_auto_node_in_in_a_bits_data; 
  wire  sbypass_auto_node_in_in_a_bits_corrupt; 
  wire  sbypass_auto_node_in_in_d_ready; 
  wire  sbypass_auto_node_in_in_d_valid; 
  wire [2:0] sbypass_auto_node_in_in_d_bits_opcode; 
  wire [1:0] sbypass_auto_node_in_in_d_bits_param; 
  wire [2:0] sbypass_auto_node_in_in_d_bits_size; 
  wire [2:0] sbypass_auto_node_in_in_d_bits_source; 
  wire [4:0] sbypass_auto_node_in_in_d_bits_sink; 
  wire  sbypass_auto_node_in_in_d_bits_denied; 
  wire [31:0] sbypass_auto_node_in_in_d_bits_data; 
  wire  sbypass_auto_node_in_in_d_bits_corrupt; 
  wire  sbypass_io_bypass; 
  wire  mbypass_clock; 
  wire  mbypass_reset; 
  wire  mbypass_auto_in_1_a_ready; 
  wire  mbypass_auto_in_1_a_valid; 
  wire [2:0] mbypass_auto_in_1_a_bits_opcode; 
  wire [2:0] mbypass_auto_in_1_a_bits_param; 
  wire [3:0] mbypass_auto_in_1_a_bits_size; 
  wire [5:0] mbypass_auto_in_1_a_bits_source; 
  wire [31:0] mbypass_auto_in_1_a_bits_address; 
  wire [3:0] mbypass_auto_in_1_a_bits_mask; 
  wire [31:0] mbypass_auto_in_1_a_bits_data; 
  wire  mbypass_auto_in_1_c_ready; 
  wire  mbypass_auto_in_1_c_valid; 
  wire [2:0] mbypass_auto_in_1_c_bits_opcode; 
  wire [2:0] mbypass_auto_in_1_c_bits_param; 
  wire [3:0] mbypass_auto_in_1_c_bits_size; 
  wire [5:0] mbypass_auto_in_1_c_bits_source; 
  wire [31:0] mbypass_auto_in_1_c_bits_address; 
  wire  mbypass_auto_in_1_d_ready; 
  wire  mbypass_auto_in_1_d_valid; 
  wire [2:0] mbypass_auto_in_1_d_bits_opcode; 
  wire [1:0] mbypass_auto_in_1_d_bits_param; 
  wire [3:0] mbypass_auto_in_1_d_bits_size; 
  wire [5:0] mbypass_auto_in_1_d_bits_source; 
  wire  mbypass_auto_in_1_d_bits_sink; 
  wire  mbypass_auto_in_1_d_bits_denied; 
  wire [31:0] mbypass_auto_in_1_d_bits_data; 
  wire  mbypass_auto_in_1_e_ready; 
  wire  mbypass_auto_in_1_e_valid; 
  wire  mbypass_auto_in_1_e_bits_sink; 
  wire  mbypass_auto_in_0_c_ready; 
  wire  mbypass_auto_in_0_c_valid; 
  wire [2:0] mbypass_auto_in_0_c_bits_opcode; 
  wire [2:0] mbypass_auto_in_0_c_bits_param; 
  wire [3:0] mbypass_auto_in_0_c_bits_size; 
  wire  mbypass_auto_in_0_c_bits_source; 
  wire [31:0] mbypass_auto_in_0_c_bits_address; 
  wire  mbypass_auto_in_0_c_bits_corrupt; 
  wire  mbypass_auto_in_0_d_valid; 
  wire [2:0] mbypass_auto_in_0_d_bits_opcode; 
  wire [1:0] mbypass_auto_in_0_d_bits_param; 
  wire [3:0] mbypass_auto_in_0_d_bits_size; 
  wire  mbypass_auto_in_0_d_bits_source; 
  wire  mbypass_auto_in_0_d_bits_sink; 
  wire  mbypass_auto_in_0_d_bits_denied; 
  wire  mbypass_auto_in_0_d_bits_corrupt; 
  wire  mbypass_auto_out_a_ready; 
  wire  mbypass_auto_out_a_valid; 
  wire [2:0] mbypass_auto_out_a_bits_opcode; 
  wire [2:0] mbypass_auto_out_a_bits_param; 
  wire [3:0] mbypass_auto_out_a_bits_size; 
  wire [5:0] mbypass_auto_out_a_bits_source; 
  wire [31:0] mbypass_auto_out_a_bits_address; 
  wire [3:0] mbypass_auto_out_a_bits_mask; 
  wire [31:0] mbypass_auto_out_a_bits_data; 
  wire  mbypass_auto_out_c_ready; 
  wire  mbypass_auto_out_c_valid; 
  wire [2:0] mbypass_auto_out_c_bits_opcode; 
  wire [2:0] mbypass_auto_out_c_bits_param; 
  wire [3:0] mbypass_auto_out_c_bits_size; 
  wire [5:0] mbypass_auto_out_c_bits_source; 
  wire [31:0] mbypass_auto_out_c_bits_address; 
  wire  mbypass_auto_out_c_bits_corrupt; 
  wire  mbypass_auto_out_d_ready; 
  wire  mbypass_auto_out_d_valid; 
  wire [2:0] mbypass_auto_out_d_bits_opcode; 
  wire [1:0] mbypass_auto_out_d_bits_param; 
  wire [3:0] mbypass_auto_out_d_bits_size; 
  wire [5:0] mbypass_auto_out_d_bits_source; 
  wire  mbypass_auto_out_d_bits_sink; 
  wire  mbypass_auto_out_d_bits_denied; 
  wire [31:0] mbypass_auto_out_d_bits_data; 
  wire  mbypass_auto_out_d_bits_corrupt; 
  wire  mbypass_auto_out_e_ready; 
  wire  mbypass_auto_out_e_valid; 
  wire  mbypass_auto_out_e_bits_sink; 
  wire  mbypass_io_bypass; 
  wire  buffer_clock; 
  wire  buffer_reset; 
  wire  buffer_auto_out_c_ready; 
  wire  buffer_auto_out_c_valid; 
  wire [2:0] buffer_auto_out_c_bits_opcode; 
  wire [2:0] buffer_auto_out_c_bits_param; 
  wire [3:0] buffer_auto_out_c_bits_size; 
  wire  buffer_auto_out_c_bits_source; 
  wire [31:0] buffer_auto_out_c_bits_address; 
  wire  buffer_auto_out_c_bits_corrupt; 
  wire  buffer_auto_out_d_valid; 
  wire [2:0] buffer_auto_out_d_bits_opcode; 
  wire [1:0] buffer_auto_out_d_bits_param; 
  wire [3:0] buffer_auto_out_d_bits_size; 
  wire  buffer_auto_out_d_bits_source; 
  wire  buffer_auto_out_d_bits_sink; 
  wire  buffer_auto_out_d_bits_denied; 
  wire  buffer_auto_out_d_bits_corrupt; 
  wire  TLMonitor_clock; 
  wire  TLMonitor_reset; 
  wire  TLMonitor_io_in_a_ready; 
  wire  TLMonitor_io_in_a_valid; 
  wire [2:0] TLMonitor_io_in_a_bits_opcode; 
  wire [2:0] TLMonitor_io_in_a_bits_param; 
  wire [2:0] TLMonitor_io_in_a_bits_size; 
  wire [2:0] TLMonitor_io_in_a_bits_source; 
  wire [31:0] TLMonitor_io_in_a_bits_address; 
  wire [3:0] TLMonitor_io_in_a_bits_mask; 
  wire  TLMonitor_io_in_a_bits_corrupt; 
  wire  TLMonitor_io_in_bvalid; 
  wire  TLMonitor_io_in_d_ready; 
  wire  TLMonitor_io_in_d_valid; 
  wire [2:0] TLMonitor_io_in_d_bits_opcode; 
  wire [1:0] TLMonitor_io_in_d_bits_param; 
  wire [2:0] TLMonitor_io_in_d_bits_size; 
  wire [2:0] TLMonitor_io_in_d_bits_source; 
  wire [4:0] TLMonitor_io_in_d_bits_sink; 
  wire  TLMonitor_io_in_d_bits_denied; 
  wire  TLMonitor_io_in_d_bits_corrupt; 
  wire  sinkA_clock; 
  wire  sinkA_reset; 
  wire  sinkA_io_a_ready; 
  wire  sinkA_io_a_valid; 
  wire [2:0] sinkA_io_a_bits_opcode; 
  wire [2:0] sinkA_io_a_bits_param; 
  wire [2:0] sinkA_io_a_bits_size; 
  wire [2:0] sinkA_io_a_bits_source; 
  wire [31:0] sinkA_io_a_bits_address; 
  wire [3:0] sinkA_io_a_bits_mask; 
  wire [31:0] sinkA_io_a_bits_data; 
  wire  sinkA_io_q_ready; 
  wire  sinkA_io_q_valid; 
  wire [31:0] sinkA_io_q_bits_data; 
  wire  sinkA_io_q_bits_last; 
  wire [12:0] sinkA_io_q_bits_beats; 
  wire  sinkB_clock; 
  wire  sinkB_reset; 
  wire  sinkB_io_q_ready; 
  wire  sinkB_io_q_valid; 
  wire [31:0] sinkB_io_q_bits_data; 
  wire  sinkB_io_q_bits_last; 
  wire  sinkC_clock; 
  wire  sinkC_reset; 
  wire  sinkC_io_q_ready; 
  wire  sinkC_io_q_valid; 
  wire [31:0] sinkC_io_q_bits_data; 
  wire  sinkC_io_q_bits_last; 
  wire  sinkD_clock; 
  wire  sinkD_reset; 
  wire  sinkD_io_d_ready; 
  wire  sinkD_io_d_valid; 
  wire [2:0] sinkD_io_d_bits_opcode; 
  wire [1:0] sinkD_io_d_bits_param; 
  wire [3:0] sinkD_io_d_bits_size; 
  wire [5:0] sinkD_io_d_bits_source; 
  wire  sinkD_io_d_bits_sink; 
  wire  sinkD_io_d_bits_denied; 
  wire [31:0] sinkD_io_d_bits_data; 
  wire  sinkD_io_q_ready; 
  wire  sinkD_io_q_valid; 
  wire [31:0] sinkD_io_q_bits_data; 
  wire  sinkD_io_q_bits_last; 
  wire [12:0] sinkD_io_q_bits_beats; 
  wire  sinkD_io_a_tlSource_valid; 
  wire [5:0] sinkD_io_a_tlSource_bits; 
  wire [15:0] sinkD_io_a_clSource; 
  wire  sinkD_io_c_tlSource_valid; 
  wire [5:0] sinkD_io_c_tlSource_bits; 
  wire [15:0] sinkD_io_c_clSource; 
  wire [31:0] sinkE_io_q_bits_data; 
  wire [15:0] sinkE_io_d_clSink; 
  wire  sourceA_clock; 
  wire  sourceA_reset; 
  wire  sourceA_io_a_ready; 
  wire  sourceA_io_a_valid; 
  wire [2:0] sourceA_io_a_bits_opcode; 
  wire [2:0] sourceA_io_a_bits_param; 
  wire [3:0] sourceA_io_a_bits_size; 
  wire [5:0] sourceA_io_a_bits_source; 
  wire [31:0] sourceA_io_a_bits_address; 
  wire [3:0] sourceA_io_a_bits_mask; 
  wire [31:0] sourceA_io_a_bits_data; 
  wire  sourceA_io_q_ready; 
  wire  sourceA_io_q_valid; 
  wire [31:0] sourceA_io_q_bits; 
  wire  sourceA_io_d_tlSource_valid; 
  wire [5:0] sourceA_io_d_tlSource_bits; 
  wire [15:0] sourceA_io_d_clSource; 
  wire  sourceB_clock; 
  wire  sourceB_reset; 
  wire  sourceB_io_bvalid; 
  wire  sourceB_io_q_ready; 
  wire  sourceB_io_q_valid; 
  wire [31:0] sourceB_io_q_bits; 
  wire  sourceC_clock; 
  wire  sourceC_reset; 
  wire  sourceC_io_c_ready; 
  wire  sourceC_io_c_valid; 
  wire [2:0] sourceC_io_c_bits_opcode; 
  wire [2:0] sourceC_io_c_bits_param; 
  wire [3:0] sourceC_io_c_bits_size; 
  wire [5:0] sourceC_io_c_bits_source; 
  wire [31:0] sourceC_io_c_bits_address; 
  wire  sourceC_io_q_ready; 
  wire  sourceC_io_q_valid; 
  wire [31:0] sourceC_io_q_bits; 
  wire  sourceC_io_d_tlSource_valid; 
  wire [5:0] sourceC_io_d_tlSource_bits; 
  wire [15:0] sourceC_io_d_clSource; 
  wire  sourceD_clock; 
  wire  sourceD_reset; 
  wire  sourceD_io_d_ready; 
  wire  sourceD_io_d_valid; 
  wire [2:0] sourceD_io_d_bits_opcode; 
  wire [1:0] sourceD_io_d_bits_param; 
  wire [2:0] sourceD_io_d_bits_size; 
  wire [2:0] sourceD_io_d_bits_source; 
  wire [4:0] sourceD_io_d_bits_sink; 
  wire  sourceD_io_d_bits_denied; 
  wire [31:0] sourceD_io_d_bits_data; 
  wire  sourceD_io_d_bits_corrupt; 
  wire  sourceD_io_q_ready; 
  wire  sourceD_io_q_valid; 
  wire [31:0] sourceD_io_q_bits; 
  wire [15:0] sourceD_io_e_clSink; 
  wire  sourceE_io_e_ready; 
  wire  sourceE_io_e_valid; 
  wire  sourceE_io_e_bits_sink; 
  wire  sourceE_io_q_ready; 
  wire  sourceE_io_q_valid; 
  wire [31:0] sourceE_io_q_bits; 
  wire  rx_clock; 
  wire  rx_reset; 
  wire  rx_io_b2c_send; 
  wire [31:0] rx_io_b2c_data; 
  wire [31:0] rx_io_a_mem_0; 
  wire [31:0] rx_io_a_mem_1; 
  wire [31:0] rx_io_a_mem_2; 
  wire [31:0] rx_io_a_mem_3; 
  wire [31:0] rx_io_a_mem_4; 
  wire [31:0] rx_io_a_mem_5; 
  wire [31:0] rx_io_a_mem_6; 
  wire [31:0] rx_io_a_mem_7; 
  wire [3:0] rx_io_a_ridx; 
  wire [3:0] rx_io_a_widx; 
  wire  rx_io_a_safe_ridx_valid; 
  wire  rx_io_a_safe_widx_valid; 
  wire  rx_io_a_safe_source_reset_n; 
  wire  rx_io_a_safe_sink_reset_n; 
  wire [31:0] rx_io_bmem_0; 
  wire [31:0] rx_io_bmem_1; 
  wire [31:0] rx_io_bmem_2; 
  wire [31:0] rx_io_bmem_3; 
  wire [31:0] rx_io_bmem_4; 
  wire [31:0] rx_io_bmem_5; 
  wire [31:0] rx_io_bmem_6; 
  wire [31:0] rx_io_bmem_7; 
  wire [3:0] rx_io_bridx; 
  wire [3:0] rx_io_bwidx; 
  wire  rx_io_bsafe_ridx_valid; 
  wire  rx_io_bsafe_widx_valid; 
  wire  rx_io_bsafe_source_reset_n; 
  wire  rx_io_bsafe_sink_reset_n; 
  wire [31:0] rx_io_c_mem_0; 
  wire [31:0] rx_io_c_mem_1; 
  wire [31:0] rx_io_c_mem_2; 
  wire [31:0] rx_io_c_mem_3; 
  wire [31:0] rx_io_c_mem_4; 
  wire [31:0] rx_io_c_mem_5; 
  wire [31:0] rx_io_c_mem_6; 
  wire [31:0] rx_io_c_mem_7; 
  wire [3:0] rx_io_c_ridx; 
  wire [3:0] rx_io_c_widx; 
  wire  rx_io_c_safe_ridx_valid; 
  wire  rx_io_c_safe_widx_valid; 
  wire  rx_io_c_safe_source_reset_n; 
  wire  rx_io_c_safe_sink_reset_n; 
  wire [31:0] rx_io_d_mem_0; 
  wire [31:0] rx_io_d_mem_1; 
  wire [31:0] rx_io_d_mem_2; 
  wire [31:0] rx_io_d_mem_3; 
  wire [31:0] rx_io_d_mem_4; 
  wire [31:0] rx_io_d_mem_5; 
  wire [31:0] rx_io_d_mem_6; 
  wire [31:0] rx_io_d_mem_7; 
  wire [3:0] rx_io_d_ridx; 
  wire [3:0] rx_io_d_widx; 
  wire  rx_io_d_safe_ridx_valid; 
  wire  rx_io_d_safe_widx_valid; 
  wire  rx_io_d_safe_source_reset_n; 
  wire  rx_io_d_safe_sink_reset_n; 
  wire [31:0] rx_io_e_mem_0; 
  wire [31:0] rx_io_e_mem_1; 
  wire [31:0] rx_io_e_mem_2; 
  wire [31:0] rx_io_e_mem_3; 
  wire [31:0] rx_io_e_mem_4; 
  wire [31:0] rx_io_e_mem_5; 
  wire [31:0] rx_io_e_mem_6; 
  wire [31:0] rx_io_e_mem_7; 
  wire [3:0] rx_io_e_ridx; 
  wire [3:0] rx_io_e_widx; 
  wire  rx_io_e_safe_ridx_valid; 
  wire  rx_io_e_safe_widx_valid; 
  wire  rx_io_e_safe_source_reset_n; 
  wire  rx_io_e_safe_sink_reset_n; 
  wire [19:0] rx_io_rxc_mem_0_a; 
  wire [19:0] rx_io_rxc_mem_0_b; 
  wire [19:0] rx_io_rxc_mem_0_c; 
  wire [19:0] rx_io_rxc_mem_0_d; 
  wire [19:0] rx_io_rxc_mem_0_e; 
  wire  rx_io_rxc_ridx; 
  wire  rx_io_rxc_widx; 
  wire  rx_io_rxc_safe_ridx_valid; 
  wire  rx_io_rxc_safe_widx_valid; 
  wire  rx_io_rxc_safe_source_reset_n; 
  wire  rx_io_rxc_safe_sink_reset_n; 
  wire [19:0] rx_io_txc_mem_0_a; 
  wire [19:0] rx_io_txc_mem_0_b; 
  wire [19:0] rx_io_txc_mem_0_c; 
  wire [19:0] rx_io_txc_mem_0_d; 
  wire [19:0] rx_io_txc_mem_0_e; 
  wire  rx_io_txc_ridx; 
  wire  rx_io_txc_widx; 
  wire  rx_io_txc_safe_ridx_valid; 
  wire  rx_io_txc_safe_widx_valid; 
  wire  rx_io_txc_safe_source_reset_n; 
  wire  rx_io_txc_safe_sink_reset_n; 
  wire  AsyncResetReg_d; 
  wire  AsyncResetReg_q; 
  wire  AsyncResetReg_en; 
  wire  AsyncResetReg_clk; 
  wire  AsyncResetReg_rst; 
  wire  AsyncQueueSink_clock; 
  wire  AsyncQueueSink_reset; 
  wire  AsyncQueueSink_io_deq_ready; 
  wire  AsyncQueueSink_io_deq_valid; 
  wire [31:0] AsyncQueueSink_io_deq_bits; 
  wire [31:0] AsyncQueueSink_io_async_mem_0; 
  wire [31:0] AsyncQueueSink_io_async_mem_1; 
  wire [31:0] AsyncQueueSink_io_async_mem_2; 
  wire [31:0] AsyncQueueSink_io_async_mem_3; 
  wire [31:0] AsyncQueueSink_io_async_mem_4; 
  wire [31:0] AsyncQueueSink_io_async_mem_5; 
  wire [31:0] AsyncQueueSink_io_async_mem_6; 
  wire [31:0] AsyncQueueSink_io_async_mem_7; 
  wire [3:0] AsyncQueueSink_io_async_ridx; 
  wire [3:0] AsyncQueueSink_io_async_widx; 
  wire  AsyncQueueSink_io_async_safe_ridx_valid; 
  wire  AsyncQueueSink_io_async_safe_widx_valid; 
  wire  AsyncQueueSink_io_async_safe_source_reset_n; 
  wire  AsyncQueueSink_io_async_safe_sink_reset_n; 
  wire  AsyncQueueSink_1_clock; 
  wire  AsyncQueueSink_1_reset; 
  wire  AsyncQueueSink_1_io_deq_ready; 
  wire  AsyncQueueSink_1_io_deq_valid; 
  wire [31:0] AsyncQueueSink_1_io_deq_bits; 
  wire [31:0] AsyncQueueSink_1_io_async_mem_0; 
  wire [31:0] AsyncQueueSink_1_io_async_mem_1; 
  wire [31:0] AsyncQueueSink_1_io_async_mem_2; 
  wire [31:0] AsyncQueueSink_1_io_async_mem_3; 
  wire [31:0] AsyncQueueSink_1_io_async_mem_4; 
  wire [31:0] AsyncQueueSink_1_io_async_mem_5; 
  wire [31:0] AsyncQueueSink_1_io_async_mem_6; 
  wire [31:0] AsyncQueueSink_1_io_async_mem_7; 
  wire [3:0] AsyncQueueSink_1_io_async_ridx; 
  wire [3:0] AsyncQueueSink_1_io_async_widx; 
  wire  AsyncQueueSink_1_io_async_safe_ridx_valid; 
  wire  AsyncQueueSink_1_io_async_safe_widx_valid; 
  wire  AsyncQueueSink_1_io_async_safe_source_reset_n; 
  wire  AsyncQueueSink_1_io_async_safe_sink_reset_n; 
  wire  AsyncQueueSink_2_clock; 
  wire  AsyncQueueSink_2_reset; 
  wire  AsyncQueueSink_2_io_deq_ready; 
  wire  AsyncQueueSink_2_io_deq_valid; 
  wire [31:0] AsyncQueueSink_2_io_deq_bits; 
  wire [31:0] AsyncQueueSink_2_io_async_mem_0; 
  wire [31:0] AsyncQueueSink_2_io_async_mem_1; 
  wire [31:0] AsyncQueueSink_2_io_async_mem_2; 
  wire [31:0] AsyncQueueSink_2_io_async_mem_3; 
  wire [31:0] AsyncQueueSink_2_io_async_mem_4; 
  wire [31:0] AsyncQueueSink_2_io_async_mem_5; 
  wire [31:0] AsyncQueueSink_2_io_async_mem_6; 
  wire [31:0] AsyncQueueSink_2_io_async_mem_7; 
  wire [3:0] AsyncQueueSink_2_io_async_ridx; 
  wire [3:0] AsyncQueueSink_2_io_async_widx; 
  wire  AsyncQueueSink_2_io_async_safe_ridx_valid; 
  wire  AsyncQueueSink_2_io_async_safe_widx_valid; 
  wire  AsyncQueueSink_2_io_async_safe_source_reset_n; 
  wire  AsyncQueueSink_2_io_async_safe_sink_reset_n; 
  wire  AsyncQueueSink_3_clock; 
  wire  AsyncQueueSink_3_reset; 
  wire  AsyncQueueSink_3_io_deq_ready; 
  wire  AsyncQueueSink_3_io_deq_valid; 
  wire [31:0] AsyncQueueSink_3_io_deq_bits; 
  wire [31:0] AsyncQueueSink_3_io_async_mem_0; 
  wire [31:0] AsyncQueueSink_3_io_async_mem_1; 
  wire [31:0] AsyncQueueSink_3_io_async_mem_2; 
  wire [31:0] AsyncQueueSink_3_io_async_mem_3; 
  wire [31:0] AsyncQueueSink_3_io_async_mem_4; 
  wire [31:0] AsyncQueueSink_3_io_async_mem_5; 
  wire [31:0] AsyncQueueSink_3_io_async_mem_6; 
  wire [31:0] AsyncQueueSink_3_io_async_mem_7; 
  wire [3:0] AsyncQueueSink_3_io_async_ridx; 
  wire [3:0] AsyncQueueSink_3_io_async_widx; 
  wire  AsyncQueueSink_3_io_async_safe_ridx_valid; 
  wire  AsyncQueueSink_3_io_async_safe_widx_valid; 
  wire  AsyncQueueSink_3_io_async_safe_source_reset_n; 
  wire  AsyncQueueSink_3_io_async_safe_sink_reset_n; 
  wire  AsyncQueueSink_4_clock; 
  wire  AsyncQueueSink_4_reset; 
  wire  AsyncQueueSink_4_io_deq_ready; 
  wire  AsyncQueueSink_4_io_deq_valid; 
  wire [31:0] AsyncQueueSink_4_io_deq_bits; 
  wire [31:0] AsyncQueueSink_4_io_async_mem_0; 
  wire [31:0] AsyncQueueSink_4_io_async_mem_1; 
  wire [31:0] AsyncQueueSink_4_io_async_mem_2; 
  wire [31:0] AsyncQueueSink_4_io_async_mem_3; 
  wire [31:0] AsyncQueueSink_4_io_async_mem_4; 
  wire [31:0] AsyncQueueSink_4_io_async_mem_5; 
  wire [31:0] AsyncQueueSink_4_io_async_mem_6; 
  wire [31:0] AsyncQueueSink_4_io_async_mem_7; 
  wire [3:0] AsyncQueueSink_4_io_async_ridx; 
  wire [3:0] AsyncQueueSink_4_io_async_widx; 
  wire  AsyncQueueSink_4_io_async_safe_ridx_valid; 
  wire  AsyncQueueSink_4_io_async_safe_widx_valid; 
  wire  AsyncQueueSink_4_io_async_safe_source_reset_n; 
  wire  AsyncQueueSink_4_io_async_safe_sink_reset_n; 
  wire  tx_clock; 
  wire  tx_reset; 
  wire  tx_io_c2b_clk; 
  wire  tx_io_c2b_rst; 
  wire  tx_io_c2b_send; 
  wire [31:0] tx_io_c2b_data; 
  wire  tx_io_sa_ready; 
  wire  tx_io_sa_valid; 
  wire [31:0] tx_io_sa_bits_data; 
  wire  tx_io_sa_bits_last; 
  wire [12:0] tx_io_sa_bits_beats; 
  wire  tx_io_sb_ready; 
  wire [31:0] tx_io_sb_bits_data; 
  wire  tx_io_sb_bits_last; 
  wire  tx_io_sc_ready; 
  wire [31:0] tx_io_sc_bits_data; 
  wire  tx_io_sc_bits_last; 
  wire  tx_io_sd_ready; 
  wire  tx_io_sd_valid; 
  wire [31:0] tx_io_sd_bits_data; 
  wire  tx_io_sd_bits_last; 
  wire [12:0] tx_io_sd_bits_beats; 
  wire [31:0] tx_io_se_bits_data; 
  wire [19:0] tx_io_rxc_mem_0_a; 
  wire [19:0] tx_io_rxc_mem_0_b; 
  wire [19:0] tx_io_rxc_mem_0_c; 
  wire [19:0] tx_io_rxc_mem_0_d; 
  wire [19:0] tx_io_rxc_mem_0_e; 
  wire  tx_io_rxc_ridx; 
  wire  tx_io_rxc_widx; 
  wire  tx_io_rxc_safe_ridx_valid; 
  wire  tx_io_rxc_safe_widx_valid; 
  wire  tx_io_rxc_safe_source_reset_n; 
  wire  tx_io_rxc_safe_sink_reset_n; 
  wire [19:0] tx_io_txc_mem_0_a; 
  wire [19:0] tx_io_txc_mem_0_b; 
  wire [19:0] tx_io_txc_mem_0_c; 
  wire [19:0] tx_io_txc_mem_0_d; 
  wire [19:0] tx_io_txc_mem_0_e; 
  wire  tx_io_txc_ridx; 
  wire  tx_io_txc_widx; 
  wire  tx_io_txc_safe_ridx_valid; 
  wire  tx_io_txc_safe_widx_valid; 
  wire  tx_io_txc_safe_source_reset_n; 
  wire  tx_io_txc_safe_sink_reset_n; 
  wire  ResetCatchAndSync_d3_clock; 
  wire  ResetCatchAndSync_d3_reset; 
  wire  ResetCatchAndSync_d3_io_sync_reset; 
  wire  ResetCatchAndSync_d3_1_clock; 
  wire  ResetCatchAndSync_d3_1_reset; 
  wire  ResetCatchAndSync_d3_1_io_sync_reset; 
  dual_TLBusBypass sbypass ( 
    .clock(sbypass_clock),
    .reset(sbypass_reset),
    .auto_node_out_out_a_ready(sbypass_auto_node_out_out_a_ready),
    .auto_node_out_out_a_valid(sbypass_auto_node_out_out_a_valid),
    .auto_node_out_out_a_bits_opcode(sbypass_auto_node_out_out_a_bits_opcode),
    .auto_node_out_out_a_bits_param(sbypass_auto_node_out_out_a_bits_param),
    .auto_node_out_out_a_bits_size(sbypass_auto_node_out_out_a_bits_size),
    .auto_node_out_out_a_bits_source(sbypass_auto_node_out_out_a_bits_source),
    .auto_node_out_out_a_bits_address(sbypass_auto_node_out_out_a_bits_address),
    .auto_node_out_out_a_bits_mask(sbypass_auto_node_out_out_a_bits_mask),
    .auto_node_out_out_a_bits_data(sbypass_auto_node_out_out_a_bits_data),
    .auto_node_out_out_a_bits_corrupt(sbypass_auto_node_out_out_a_bits_corrupt),
    .auto_node_out_out_d_ready(sbypass_auto_node_out_out_d_ready),
    .auto_node_out_out_d_valid(sbypass_auto_node_out_out_d_valid),
    .auto_node_out_out_d_bits_opcode(sbypass_auto_node_out_out_d_bits_opcode),
    .auto_node_out_out_d_bits_param(sbypass_auto_node_out_out_d_bits_param),
    .auto_node_out_out_d_bits_size(sbypass_auto_node_out_out_d_bits_size),
    .auto_node_out_out_d_bits_source(sbypass_auto_node_out_out_d_bits_source),
    .auto_node_out_out_d_bits_sink(sbypass_auto_node_out_out_d_bits_sink),
    .auto_node_out_out_d_bits_denied(sbypass_auto_node_out_out_d_bits_denied),
    .auto_node_out_out_d_bits_data(sbypass_auto_node_out_out_d_bits_data),
    .auto_node_out_out_d_bits_corrupt(sbypass_auto_node_out_out_d_bits_corrupt),
    .auto_node_in_in_a_ready(sbypass_auto_node_in_in_a_ready),
    .auto_node_in_in_a_valid(sbypass_auto_node_in_in_a_valid),
    .auto_node_in_in_a_bits_opcode(sbypass_auto_node_in_in_a_bits_opcode),
    .auto_node_in_in_a_bits_param(sbypass_auto_node_in_in_a_bits_param),
    .auto_node_in_in_a_bits_size(sbypass_auto_node_in_in_a_bits_size),
    .auto_node_in_in_a_bits_source(sbypass_auto_node_in_in_a_bits_source),
    .auto_node_in_in_a_bits_address(sbypass_auto_node_in_in_a_bits_address),
    .auto_node_in_in_a_bits_mask(sbypass_auto_node_in_in_a_bits_mask),
    .auto_node_in_in_a_bits_data(sbypass_auto_node_in_in_a_bits_data),
    .auto_node_in_in_a_bits_corrupt(sbypass_auto_node_in_in_a_bits_corrupt),
    .auto_node_in_in_d_ready(sbypass_auto_node_in_in_d_ready),
    .auto_node_in_in_d_valid(sbypass_auto_node_in_in_d_valid),
    .auto_node_in_in_d_bits_opcode(sbypass_auto_node_in_in_d_bits_opcode),
    .auto_node_in_in_d_bits_param(sbypass_auto_node_in_in_d_bits_param),
    .auto_node_in_in_d_bits_size(sbypass_auto_node_in_in_d_bits_size),
    .auto_node_in_in_d_bits_source(sbypass_auto_node_in_in_d_bits_source),
    .auto_node_in_in_d_bits_sink(sbypass_auto_node_in_in_d_bits_sink),
    .auto_node_in_in_d_bits_denied(sbypass_auto_node_in_in_d_bits_denied),
    .auto_node_in_in_d_bits_data(sbypass_auto_node_in_in_d_bits_data),
    .auto_node_in_in_d_bits_corrupt(sbypass_auto_node_in_in_d_bits_corrupt),
    .io_bypass(sbypass_io_bypass)
  );
  dual_MasterMux mbypass ( 
    .clock(mbypass_clock),
    .reset(mbypass_reset),
    .auto_in_1_a_ready(mbypass_auto_in_1_a_ready),
    .auto_in_1_a_valid(mbypass_auto_in_1_a_valid),
    .auto_in_1_a_bits_opcode(mbypass_auto_in_1_a_bits_opcode),
    .auto_in_1_a_bits_param(mbypass_auto_in_1_a_bits_param),
    .auto_in_1_a_bits_size(mbypass_auto_in_1_a_bits_size),
    .auto_in_1_a_bits_source(mbypass_auto_in_1_a_bits_source),
    .auto_in_1_a_bits_address(mbypass_auto_in_1_a_bits_address),
    .auto_in_1_a_bits_mask(mbypass_auto_in_1_a_bits_mask),
    .auto_in_1_a_bits_data(mbypass_auto_in_1_a_bits_data),
    .auto_in_1_c_ready(mbypass_auto_in_1_c_ready),
    .auto_in_1_c_valid(mbypass_auto_in_1_c_valid),
    .auto_in_1_c_bits_opcode(mbypass_auto_in_1_c_bits_opcode),
    .auto_in_1_c_bits_param(mbypass_auto_in_1_c_bits_param),
    .auto_in_1_c_bits_size(mbypass_auto_in_1_c_bits_size),
    .auto_in_1_c_bits_source(mbypass_auto_in_1_c_bits_source),
    .auto_in_1_c_bits_address(mbypass_auto_in_1_c_bits_address),
    .auto_in_1_d_ready(mbypass_auto_in_1_d_ready),
    .auto_in_1_d_valid(mbypass_auto_in_1_d_valid),
    .auto_in_1_d_bits_opcode(mbypass_auto_in_1_d_bits_opcode),
    .auto_in_1_d_bits_param(mbypass_auto_in_1_d_bits_param),
    .auto_in_1_d_bits_size(mbypass_auto_in_1_d_bits_size),
    .auto_in_1_d_bits_source(mbypass_auto_in_1_d_bits_source),
    .auto_in_1_d_bits_sink(mbypass_auto_in_1_d_bits_sink),
    .auto_in_1_d_bits_denied(mbypass_auto_in_1_d_bits_denied),
    .auto_in_1_d_bits_data(mbypass_auto_in_1_d_bits_data),
    .auto_in_1_e_ready(mbypass_auto_in_1_e_ready),
    .auto_in_1_e_valid(mbypass_auto_in_1_e_valid),
    .auto_in_1_e_bits_sink(mbypass_auto_in_1_e_bits_sink),
    .auto_in_0_c_ready(mbypass_auto_in_0_c_ready),
    .auto_in_0_c_valid(mbypass_auto_in_0_c_valid),
    .auto_in_0_c_bits_opcode(mbypass_auto_in_0_c_bits_opcode),
    .auto_in_0_c_bits_param(mbypass_auto_in_0_c_bits_param),
    .auto_in_0_c_bits_size(mbypass_auto_in_0_c_bits_size),
    .auto_in_0_c_bits_source(mbypass_auto_in_0_c_bits_source),
    .auto_in_0_c_bits_address(mbypass_auto_in_0_c_bits_address),
    .auto_in_0_c_bits_corrupt(mbypass_auto_in_0_c_bits_corrupt),
    .auto_in_0_d_valid(mbypass_auto_in_0_d_valid),
    .auto_in_0_d_bits_opcode(mbypass_auto_in_0_d_bits_opcode),
    .auto_in_0_d_bits_param(mbypass_auto_in_0_d_bits_param),
    .auto_in_0_d_bits_size(mbypass_auto_in_0_d_bits_size),
    .auto_in_0_d_bits_source(mbypass_auto_in_0_d_bits_source),
    .auto_in_0_d_bits_sink(mbypass_auto_in_0_d_bits_sink),
    .auto_in_0_d_bits_denied(mbypass_auto_in_0_d_bits_denied),
    .auto_in_0_d_bits_corrupt(mbypass_auto_in_0_d_bits_corrupt),
    .auto_out_a_ready(mbypass_auto_out_a_ready),
    .auto_out_a_valid(mbypass_auto_out_a_valid),
    .auto_out_a_bits_opcode(mbypass_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(mbypass_auto_out_a_bits_param),
    .auto_out_a_bits_size(mbypass_auto_out_a_bits_size),
    .auto_out_a_bits_source(mbypass_auto_out_a_bits_source),
    .auto_out_a_bits_address(mbypass_auto_out_a_bits_address),
    .auto_out_a_bits_mask(mbypass_auto_out_a_bits_mask),
    .auto_out_a_bits_data(mbypass_auto_out_a_bits_data),
    .auto_out_c_ready(mbypass_auto_out_c_ready),
    .auto_out_c_valid(mbypass_auto_out_c_valid),
    .auto_out_c_bits_opcode(mbypass_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(mbypass_auto_out_c_bits_param),
    .auto_out_c_bits_size(mbypass_auto_out_c_bits_size),
    .auto_out_c_bits_source(mbypass_auto_out_c_bits_source),
    .auto_out_c_bits_address(mbypass_auto_out_c_bits_address),
    .auto_out_c_bits_corrupt(mbypass_auto_out_c_bits_corrupt),
    .auto_out_d_ready(mbypass_auto_out_d_ready),
    .auto_out_d_valid(mbypass_auto_out_d_valid),
    .auto_out_d_bits_opcode(mbypass_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(mbypass_auto_out_d_bits_param),
    .auto_out_d_bits_size(mbypass_auto_out_d_bits_size),
    .auto_out_d_bits_source(mbypass_auto_out_d_bits_source),
    .auto_out_d_bits_sink(mbypass_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(mbypass_auto_out_d_bits_denied),
    .auto_out_d_bits_data(mbypass_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(mbypass_auto_out_d_bits_corrupt),
    .auto_out_e_ready(mbypass_auto_out_e_ready),
    .auto_out_e_valid(mbypass_auto_out_e_valid),
    .auto_out_e_bits_sink(mbypass_auto_out_e_bits_sink),
    .io_bypass(mbypass_io_bypass)
  );
  dual_TLBuffer buffer ( 
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_out_c_ready(buffer_auto_out_c_ready),
    .auto_out_c_valid(buffer_auto_out_c_valid),
    .auto_out_c_bits_opcode(buffer_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(buffer_auto_out_c_bits_param),
    .auto_out_c_bits_size(buffer_auto_out_c_bits_size),
    .auto_out_c_bits_source(buffer_auto_out_c_bits_source),
    .auto_out_c_bits_address(buffer_auto_out_c_bits_address),
    .auto_out_c_bits_corrupt(buffer_auto_out_c_bits_corrupt),
    .auto_out_d_valid(buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(buffer_auto_out_d_bits_param),
    .auto_out_d_bits_size(buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_auto_out_d_bits_source),
    .auto_out_d_bits_sink(buffer_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(buffer_auto_out_d_bits_denied),
    .auto_out_d_bits_corrupt(buffer_auto_out_d_bits_corrupt)
  );
  dual_TLMonitor_8 dual_TLMonitor ( 
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_io_in_a_bits_corrupt),
    .io_in_bvalid(TLMonitor_io_in_bvalid),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt)
  );
  dual_SinkA sinkA ( 
    .clock(sinkA_clock),
    .reset(sinkA_reset),
    .io_a_ready(sinkA_io_a_ready),
    .io_a_valid(sinkA_io_a_valid),
    .io_a_bits_opcode(sinkA_io_a_bits_opcode),
    .io_a_bits_param(sinkA_io_a_bits_param),
    .io_a_bits_size(sinkA_io_a_bits_size),
    .io_a_bits_source(sinkA_io_a_bits_source),
    .io_a_bits_address(sinkA_io_a_bits_address),
    .io_a_bits_mask(sinkA_io_a_bits_mask),
    .io_a_bits_data(sinkA_io_a_bits_data),
    .io_q_ready(sinkA_io_q_ready),
    .io_q_valid(sinkA_io_q_valid),
    .io_q_bits_data(sinkA_io_q_bits_data),
    .io_q_bits_last(sinkA_io_q_bits_last),
    .io_q_bits_beats(sinkA_io_q_bits_beats)
  );
  dual_SinkB sinkB ( 
    .clock(sinkB_clock),
    .reset(sinkB_reset),
    .io_q_ready(sinkB_io_q_ready),
    .io_q_valid(sinkB_io_q_valid),
    .io_q_bits_data(sinkB_io_q_bits_data),
    .io_q_bits_last(sinkB_io_q_bits_last)
  );
  dual_SinkC sinkC ( 
    .clock(sinkC_clock),
    .reset(sinkC_reset),
    .io_q_ready(sinkC_io_q_ready),
    .io_q_valid(sinkC_io_q_valid),
    .io_q_bits_data(sinkC_io_q_bits_data),
    .io_q_bits_last(sinkC_io_q_bits_last)
  );
  dual_SinkD sinkD ( 
    .clock(sinkD_clock),
    .reset(sinkD_reset),
    .io_d_ready(sinkD_io_d_ready),
    .io_d_valid(sinkD_io_d_valid),
    .io_d_bits_opcode(sinkD_io_d_bits_opcode),
    .io_d_bits_param(sinkD_io_d_bits_param),
    .io_d_bits_size(sinkD_io_d_bits_size),
    .io_d_bits_source(sinkD_io_d_bits_source),
    .io_d_bits_sink(sinkD_io_d_bits_sink),
    .io_d_bits_denied(sinkD_io_d_bits_denied),
    .io_d_bits_data(sinkD_io_d_bits_data),
    .io_q_ready(sinkD_io_q_ready),
    .io_q_valid(sinkD_io_q_valid),
    .io_q_bits_data(sinkD_io_q_bits_data),
    .io_q_bits_last(sinkD_io_q_bits_last),
    .io_q_bits_beats(sinkD_io_q_bits_beats),
    .io_a_tlSource_valid(sinkD_io_a_tlSource_valid),
    .io_a_tlSource_bits(sinkD_io_a_tlSource_bits),
    .io_a_clSource(sinkD_io_a_clSource),
    .io_c_tlSource_valid(sinkD_io_c_tlSource_valid),
    .io_c_tlSource_bits(sinkD_io_c_tlSource_bits),
    .io_c_clSource(sinkD_io_c_clSource)
  );
  dual_SinkE sinkE ( 
    .io_q_bits_data(sinkE_io_q_bits_data),
    .io_d_clSink(sinkE_io_d_clSink)
  );
  dual_SourceA sourceA ( 
    .clock(sourceA_clock),
    .reset(sourceA_reset),
    .io_a_ready(sourceA_io_a_ready),
    .io_a_valid(sourceA_io_a_valid),
    .io_a_bits_opcode(sourceA_io_a_bits_opcode),
    .io_a_bits_param(sourceA_io_a_bits_param),
    .io_a_bits_size(sourceA_io_a_bits_size),
    .io_a_bits_source(sourceA_io_a_bits_source),
    .io_a_bits_address(sourceA_io_a_bits_address),
    .io_a_bits_mask(sourceA_io_a_bits_mask),
    .io_a_bits_data(sourceA_io_a_bits_data),
    .io_q_ready(sourceA_io_q_ready),
    .io_q_valid(sourceA_io_q_valid),
    .io_q_bits(sourceA_io_q_bits),
    .io_d_tlSource_valid(sourceA_io_d_tlSource_valid),
    .io_d_tlSource_bits(sourceA_io_d_tlSource_bits),
    .io_d_clSource(sourceA_io_d_clSource)
  );
  dual_SourceB sourceB ( 
    .clock(sourceB_clock),
    .reset(sourceB_reset),
    .io_bvalid(sourceB_io_bvalid),
    .io_q_ready(sourceB_io_q_ready),
    .io_q_valid(sourceB_io_q_valid),
    .io_q_bits(sourceB_io_q_bits)
  );
  dual_SourceC sourceC ( 
    .clock(sourceC_clock),
    .reset(sourceC_reset),
    .io_c_ready(sourceC_io_c_ready),
    .io_c_valid(sourceC_io_c_valid),
    .io_c_bits_opcode(sourceC_io_c_bits_opcode),
    .io_c_bits_param(sourceC_io_c_bits_param),
    .io_c_bits_size(sourceC_io_c_bits_size),
    .io_c_bits_source(sourceC_io_c_bits_source),
    .io_c_bits_address(sourceC_io_c_bits_address),
    .io_q_ready(sourceC_io_q_ready),
    .io_q_valid(sourceC_io_q_valid),
    .io_q_bits(sourceC_io_q_bits),
    .io_d_tlSource_valid(sourceC_io_d_tlSource_valid),
    .io_d_tlSource_bits(sourceC_io_d_tlSource_bits),
    .io_d_clSource(sourceC_io_d_clSource)
  );
  dual_SourceD sourceD ( 
    .clock(sourceD_clock),
    .reset(sourceD_reset),
    .io_d_ready(sourceD_io_d_ready),
    .io_d_valid(sourceD_io_d_valid),
    .io_d_bits_opcode(sourceD_io_d_bits_opcode),
    .io_d_bits_param(sourceD_io_d_bits_param),
    .io_d_bits_size(sourceD_io_d_bits_size),
    .io_d_bits_source(sourceD_io_d_bits_source),
    .io_d_bits_sink(sourceD_io_d_bits_sink),
    .io_d_bits_denied(sourceD_io_d_bits_denied),
    .io_d_bits_data(sourceD_io_d_bits_data),
    .io_d_bits_corrupt(sourceD_io_d_bits_corrupt),
    .io_q_ready(sourceD_io_q_ready),
    .io_q_valid(sourceD_io_q_valid),
    .io_q_bits(sourceD_io_q_bits),
    .io_e_clSink(sourceD_io_e_clSink)
  );
  dual_SourceE sourceE ( 
    .io_e_ready(sourceE_io_e_ready),
    .io_e_valid(sourceE_io_e_valid),
    .io_e_bits_sink(sourceE_io_e_bits_sink),
    .io_q_ready(sourceE_io_q_ready),
    .io_q_valid(sourceE_io_q_valid),
    .io_q_bits(sourceE_io_q_bits)
  );
  dual_RX rx ( 
    .clock(rx_clock),
    .reset(rx_reset),
    .io_b2c_send(rx_io_b2c_send),
    .io_b2c_data(rx_io_b2c_data),
    .io_a_mem_0(rx_io_a_mem_0),
    .io_a_mem_1(rx_io_a_mem_1),
    .io_a_mem_2(rx_io_a_mem_2),
    .io_a_mem_3(rx_io_a_mem_3),
    .io_a_mem_4(rx_io_a_mem_4),
    .io_a_mem_5(rx_io_a_mem_5),
    .io_a_mem_6(rx_io_a_mem_6),
    .io_a_mem_7(rx_io_a_mem_7),
    .io_a_ridx(rx_io_a_ridx),
    .io_a_widx(rx_io_a_widx),
    .io_a_safe_ridx_valid(rx_io_a_safe_ridx_valid),
    .io_a_safe_widx_valid(rx_io_a_safe_widx_valid),
    .io_a_safe_source_reset_n(rx_io_a_safe_source_reset_n),
    .io_a_safe_sink_reset_n(rx_io_a_safe_sink_reset_n),
    .io_bmem_0(rx_io_bmem_0),
    .io_bmem_1(rx_io_bmem_1),
    .io_bmem_2(rx_io_bmem_2),
    .io_bmem_3(rx_io_bmem_3),
    .io_bmem_4(rx_io_bmem_4),
    .io_bmem_5(rx_io_bmem_5),
    .io_bmem_6(rx_io_bmem_6),
    .io_bmem_7(rx_io_bmem_7),
    .io_bridx(rx_io_bridx),
    .io_bwidx(rx_io_bwidx),
    .io_bsafe_ridx_valid(rx_io_bsafe_ridx_valid),
    .io_bsafe_widx_valid(rx_io_bsafe_widx_valid),
    .io_bsafe_source_reset_n(rx_io_bsafe_source_reset_n),
    .io_bsafe_sink_reset_n(rx_io_bsafe_sink_reset_n),
    .io_c_mem_0(rx_io_c_mem_0),
    .io_c_mem_1(rx_io_c_mem_1),
    .io_c_mem_2(rx_io_c_mem_2),
    .io_c_mem_3(rx_io_c_mem_3),
    .io_c_mem_4(rx_io_c_mem_4),
    .io_c_mem_5(rx_io_c_mem_5),
    .io_c_mem_6(rx_io_c_mem_6),
    .io_c_mem_7(rx_io_c_mem_7),
    .io_c_ridx(rx_io_c_ridx),
    .io_c_widx(rx_io_c_widx),
    .io_c_safe_ridx_valid(rx_io_c_safe_ridx_valid),
    .io_c_safe_widx_valid(rx_io_c_safe_widx_valid),
    .io_c_safe_source_reset_n(rx_io_c_safe_source_reset_n),
    .io_c_safe_sink_reset_n(rx_io_c_safe_sink_reset_n),
    .io_d_mem_0(rx_io_d_mem_0),
    .io_d_mem_1(rx_io_d_mem_1),
    .io_d_mem_2(rx_io_d_mem_2),
    .io_d_mem_3(rx_io_d_mem_3),
    .io_d_mem_4(rx_io_d_mem_4),
    .io_d_mem_5(rx_io_d_mem_5),
    .io_d_mem_6(rx_io_d_mem_6),
    .io_d_mem_7(rx_io_d_mem_7),
    .io_d_ridx(rx_io_d_ridx),
    .io_d_widx(rx_io_d_widx),
    .io_d_safe_ridx_valid(rx_io_d_safe_ridx_valid),
    .io_d_safe_widx_valid(rx_io_d_safe_widx_valid),
    .io_d_safe_source_reset_n(rx_io_d_safe_source_reset_n),
    .io_d_safe_sink_reset_n(rx_io_d_safe_sink_reset_n),
    .io_e_mem_0(rx_io_e_mem_0),
    .io_e_mem_1(rx_io_e_mem_1),
    .io_e_mem_2(rx_io_e_mem_2),
    .io_e_mem_3(rx_io_e_mem_3),
    .io_e_mem_4(rx_io_e_mem_4),
    .io_e_mem_5(rx_io_e_mem_5),
    .io_e_mem_6(rx_io_e_mem_6),
    .io_e_mem_7(rx_io_e_mem_7),
    .io_e_ridx(rx_io_e_ridx),
    .io_e_widx(rx_io_e_widx),
    .io_e_safe_ridx_valid(rx_io_e_safe_ridx_valid),
    .io_e_safe_widx_valid(rx_io_e_safe_widx_valid),
    .io_e_safe_source_reset_n(rx_io_e_safe_source_reset_n),
    .io_e_safe_sink_reset_n(rx_io_e_safe_sink_reset_n),
    .io_rxc_mem_0_a(rx_io_rxc_mem_0_a),
    .io_rxc_mem_0_b(rx_io_rxc_mem_0_b),
    .io_rxc_mem_0_c(rx_io_rxc_mem_0_c),
    .io_rxc_mem_0_d(rx_io_rxc_mem_0_d),
    .io_rxc_mem_0_e(rx_io_rxc_mem_0_e),
    .io_rxc_ridx(rx_io_rxc_ridx),
    .io_rxc_widx(rx_io_rxc_widx),
    .io_rxc_safe_ridx_valid(rx_io_rxc_safe_ridx_valid),
    .io_rxc_safe_widx_valid(rx_io_rxc_safe_widx_valid),
    .io_rxc_safe_source_reset_n(rx_io_rxc_safe_source_reset_n),
    .io_rxc_safe_sink_reset_n(rx_io_rxc_safe_sink_reset_n),
    .io_txc_mem_0_a(rx_io_txc_mem_0_a),
    .io_txc_mem_0_b(rx_io_txc_mem_0_b),
    .io_txc_mem_0_c(rx_io_txc_mem_0_c),
    .io_txc_mem_0_d(rx_io_txc_mem_0_d),
    .io_txc_mem_0_e(rx_io_txc_mem_0_e),
    .io_txc_ridx(rx_io_txc_ridx),
    .io_txc_widx(rx_io_txc_widx),
    .io_txc_safe_ridx_valid(rx_io_txc_safe_ridx_valid),
    .io_txc_safe_widx_valid(rx_io_txc_safe_widx_valid),
    .io_txc_safe_source_reset_n(rx_io_txc_safe_source_reset_n),
    .io_txc_safe_sink_reset_n(rx_io_txc_safe_sink_reset_n)
  );
  dual_AsyncResetReg #(.RESET_VALUE(1)) AsyncResetReg ( 
    .d(AsyncResetReg_d),
    .q(AsyncResetReg_q),
    .en(AsyncResetReg_en),
    .clk(AsyncResetReg_clk),
    .rst(AsyncResetReg_rst)
  );
  dual_AsyncQueueSink AsyncQueueSink ( 
    .clock(AsyncQueueSink_clock),
    .reset(AsyncQueueSink_reset),
    .io_deq_ready(AsyncQueueSink_io_deq_ready),
    .io_deq_valid(AsyncQueueSink_io_deq_valid),
    .io_deq_bits(AsyncQueueSink_io_deq_bits),
    .io_async_mem_0(AsyncQueueSink_io_async_mem_0),
    .io_async_mem_1(AsyncQueueSink_io_async_mem_1),
    .io_async_mem_2(AsyncQueueSink_io_async_mem_2),
    .io_async_mem_3(AsyncQueueSink_io_async_mem_3),
    .io_async_mem_4(AsyncQueueSink_io_async_mem_4),
    .io_async_mem_5(AsyncQueueSink_io_async_mem_5),
    .io_async_mem_6(AsyncQueueSink_io_async_mem_6),
    .io_async_mem_7(AsyncQueueSink_io_async_mem_7),
    .io_async_ridx(AsyncQueueSink_io_async_ridx),
    .io_async_widx(AsyncQueueSink_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSink_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSink_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSink_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSink_io_async_safe_sink_reset_n)
  );
  dual_AsyncQueueSink AsyncQueueSink_1 ( 
    .clock(AsyncQueueSink_1_clock),
    .reset(AsyncQueueSink_1_reset),
    .io_deq_ready(AsyncQueueSink_1_io_deq_ready),
    .io_deq_valid(AsyncQueueSink_1_io_deq_valid),
    .io_deq_bits(AsyncQueueSink_1_io_deq_bits),
    .io_async_mem_0(AsyncQueueSink_1_io_async_mem_0),
    .io_async_mem_1(AsyncQueueSink_1_io_async_mem_1),
    .io_async_mem_2(AsyncQueueSink_1_io_async_mem_2),
    .io_async_mem_3(AsyncQueueSink_1_io_async_mem_3),
    .io_async_mem_4(AsyncQueueSink_1_io_async_mem_4),
    .io_async_mem_5(AsyncQueueSink_1_io_async_mem_5),
    .io_async_mem_6(AsyncQueueSink_1_io_async_mem_6),
    .io_async_mem_7(AsyncQueueSink_1_io_async_mem_7),
    .io_async_ridx(AsyncQueueSink_1_io_async_ridx),
    .io_async_widx(AsyncQueueSink_1_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSink_1_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSink_1_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSink_1_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSink_1_io_async_safe_sink_reset_n)
  );
  dual_AsyncQueueSink AsyncQueueSink_2 ( 
    .clock(AsyncQueueSink_2_clock),
    .reset(AsyncQueueSink_2_reset),
    .io_deq_ready(AsyncQueueSink_2_io_deq_ready),
    .io_deq_valid(AsyncQueueSink_2_io_deq_valid),
    .io_deq_bits(AsyncQueueSink_2_io_deq_bits),
    .io_async_mem_0(AsyncQueueSink_2_io_async_mem_0),
    .io_async_mem_1(AsyncQueueSink_2_io_async_mem_1),
    .io_async_mem_2(AsyncQueueSink_2_io_async_mem_2),
    .io_async_mem_3(AsyncQueueSink_2_io_async_mem_3),
    .io_async_mem_4(AsyncQueueSink_2_io_async_mem_4),
    .io_async_mem_5(AsyncQueueSink_2_io_async_mem_5),
    .io_async_mem_6(AsyncQueueSink_2_io_async_mem_6),
    .io_async_mem_7(AsyncQueueSink_2_io_async_mem_7),
    .io_async_ridx(AsyncQueueSink_2_io_async_ridx),
    .io_async_widx(AsyncQueueSink_2_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSink_2_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSink_2_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSink_2_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSink_2_io_async_safe_sink_reset_n)
  );
  dual_AsyncQueueSink AsyncQueueSink_3 ( 
    .clock(AsyncQueueSink_3_clock),
    .reset(AsyncQueueSink_3_reset),
    .io_deq_ready(AsyncQueueSink_3_io_deq_ready),
    .io_deq_valid(AsyncQueueSink_3_io_deq_valid),
    .io_deq_bits(AsyncQueueSink_3_io_deq_bits),
    .io_async_mem_0(AsyncQueueSink_3_io_async_mem_0),
    .io_async_mem_1(AsyncQueueSink_3_io_async_mem_1),
    .io_async_mem_2(AsyncQueueSink_3_io_async_mem_2),
    .io_async_mem_3(AsyncQueueSink_3_io_async_mem_3),
    .io_async_mem_4(AsyncQueueSink_3_io_async_mem_4),
    .io_async_mem_5(AsyncQueueSink_3_io_async_mem_5),
    .io_async_mem_6(AsyncQueueSink_3_io_async_mem_6),
    .io_async_mem_7(AsyncQueueSink_3_io_async_mem_7),
    .io_async_ridx(AsyncQueueSink_3_io_async_ridx),
    .io_async_widx(AsyncQueueSink_3_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSink_3_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSink_3_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSink_3_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSink_3_io_async_safe_sink_reset_n)
  );
  dual_AsyncQueueSink AsyncQueueSink_4 ( 
    .clock(AsyncQueueSink_4_clock),
    .reset(AsyncQueueSink_4_reset),
    .io_deq_ready(AsyncQueueSink_4_io_deq_ready),
    .io_deq_valid(AsyncQueueSink_4_io_deq_valid),
    .io_deq_bits(AsyncQueueSink_4_io_deq_bits),
    .io_async_mem_0(AsyncQueueSink_4_io_async_mem_0),
    .io_async_mem_1(AsyncQueueSink_4_io_async_mem_1),
    .io_async_mem_2(AsyncQueueSink_4_io_async_mem_2),
    .io_async_mem_3(AsyncQueueSink_4_io_async_mem_3),
    .io_async_mem_4(AsyncQueueSink_4_io_async_mem_4),
    .io_async_mem_5(AsyncQueueSink_4_io_async_mem_5),
    .io_async_mem_6(AsyncQueueSink_4_io_async_mem_6),
    .io_async_mem_7(AsyncQueueSink_4_io_async_mem_7),
    .io_async_ridx(AsyncQueueSink_4_io_async_ridx),
    .io_async_widx(AsyncQueueSink_4_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSink_4_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSink_4_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSink_4_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSink_4_io_async_safe_sink_reset_n)
  );
  dual_TX tx ( 
    .clock(tx_clock),
    .reset(tx_reset),
    .io_c2b_clk(tx_io_c2b_clk),
    .io_c2b_rst(tx_io_c2b_rst),
    .io_c2b_send(tx_io_c2b_send),
    .io_c2b_data(tx_io_c2b_data),
    .io_sa_ready(tx_io_sa_ready),
    .io_sa_valid(tx_io_sa_valid),
    .io_sa_bits_data(tx_io_sa_bits_data),
    .io_sa_bits_last(tx_io_sa_bits_last),
    .io_sa_bits_beats(tx_io_sa_bits_beats),
    .io_sb_ready(tx_io_sb_ready),
    .io_sb_bits_data(tx_io_sb_bits_data),
    .io_sb_bits_last(tx_io_sb_bits_last),
    .io_sc_ready(tx_io_sc_ready),
    .io_sc_bits_data(tx_io_sc_bits_data),
    .io_sc_bits_last(tx_io_sc_bits_last),
    .io_sd_ready(tx_io_sd_ready),
    .io_sd_valid(tx_io_sd_valid),
    .io_sd_bits_data(tx_io_sd_bits_data),
    .io_sd_bits_last(tx_io_sd_bits_last),
    .io_sd_bits_beats(tx_io_sd_bits_beats),
    .io_se_bits_data(tx_io_se_bits_data),
    .io_rxc_mem_0_a(tx_io_rxc_mem_0_a),
    .io_rxc_mem_0_b(tx_io_rxc_mem_0_b),
    .io_rxc_mem_0_c(tx_io_rxc_mem_0_c),
    .io_rxc_mem_0_d(tx_io_rxc_mem_0_d),
    .io_rxc_mem_0_e(tx_io_rxc_mem_0_e),
    .io_rxc_ridx(tx_io_rxc_ridx),
    .io_rxc_widx(tx_io_rxc_widx),
    .io_rxc_safe_ridx_valid(tx_io_rxc_safe_ridx_valid),
    .io_rxc_safe_widx_valid(tx_io_rxc_safe_widx_valid),
    .io_rxc_safe_source_reset_n(tx_io_rxc_safe_source_reset_n),
    .io_rxc_safe_sink_reset_n(tx_io_rxc_safe_sink_reset_n),
    .io_txc_mem_0_a(tx_io_txc_mem_0_a),
    .io_txc_mem_0_b(tx_io_txc_mem_0_b),
    .io_txc_mem_0_c(tx_io_txc_mem_0_c),
    .io_txc_mem_0_d(tx_io_txc_mem_0_d),
    .io_txc_mem_0_e(tx_io_txc_mem_0_e),
    .io_txc_ridx(tx_io_txc_ridx),
    .io_txc_widx(tx_io_txc_widx),
    .io_txc_safe_ridx_valid(tx_io_txc_safe_ridx_valid),
    .io_txc_safe_widx_valid(tx_io_txc_safe_widx_valid),
    .io_txc_safe_source_reset_n(tx_io_txc_safe_source_reset_n),
    .io_txc_safe_sink_reset_n(tx_io_txc_safe_sink_reset_n)
  );
  dual_ResetCatchAndSync_d3 ResetCatchAndSync_d3 ( 
    .clock(ResetCatchAndSync_d3_clock),
    .reset(ResetCatchAndSync_d3_reset),
    .io_sync_reset(ResetCatchAndSync_d3_io_sync_reset)
  );
  dual_ResetCatchAndSync_d3 ResetCatchAndSync_d3_1 ( 
    .clock(ResetCatchAndSync_d3_1_clock),
    .reset(ResetCatchAndSync_d3_1_reset),
    .io_sync_reset(ResetCatchAndSync_d3_1_io_sync_reset)
  );
  assign auto_mbypass_out_a_valid = mbypass_auto_out_a_valid; 
  assign auto_mbypass_out_a_bits_opcode = mbypass_auto_out_a_bits_opcode; 
  assign auto_mbypass_out_a_bits_param = mbypass_auto_out_a_bits_param; 
  assign auto_mbypass_out_a_bits_size = mbypass_auto_out_a_bits_size; 
  assign auto_mbypass_out_a_bits_source = mbypass_auto_out_a_bits_source; 
  assign auto_mbypass_out_a_bits_address = mbypass_auto_out_a_bits_address; 
  assign auto_mbypass_out_a_bits_mask = mbypass_auto_out_a_bits_mask; 
  assign auto_mbypass_out_a_bits_data = mbypass_auto_out_a_bits_data; 
  assign auto_mbypass_out_c_valid = mbypass_auto_out_c_valid; 
  assign auto_mbypass_out_c_bits_opcode = mbypass_auto_out_c_bits_opcode; 
  assign auto_mbypass_out_c_bits_param = mbypass_auto_out_c_bits_param; 
  assign auto_mbypass_out_c_bits_size = mbypass_auto_out_c_bits_size; 
  assign auto_mbypass_out_c_bits_source = mbypass_auto_out_c_bits_source; 
  assign auto_mbypass_out_c_bits_address = mbypass_auto_out_c_bits_address; 
  assign auto_mbypass_out_c_bits_corrupt = mbypass_auto_out_c_bits_corrupt; 
  assign auto_mbypass_out_d_ready = mbypass_auto_out_d_ready; 
  assign auto_mbypass_out_e_valid = mbypass_auto_out_e_valid; 
  assign auto_mbypass_out_e_bits_sink = mbypass_auto_out_e_bits_sink; 
  assign auto_sbypass_node_in_in_a_ready = sbypass_auto_node_in_in_a_ready; 
  assign auto_sbypass_node_in_in_d_valid = sbypass_auto_node_in_in_d_valid; 
  assign auto_sbypass_node_in_in_d_bits_opcode = sbypass_auto_node_in_in_d_bits_opcode; 
  assign auto_sbypass_node_in_in_d_bits_param = sbypass_auto_node_in_in_d_bits_param; 
  assign auto_sbypass_node_in_in_d_bits_size = sbypass_auto_node_in_in_d_bits_size; 
  assign auto_sbypass_node_in_in_d_bits_source = sbypass_auto_node_in_in_d_bits_source; 
  assign auto_sbypass_node_in_in_d_bits_sink = sbypass_auto_node_in_in_d_bits_sink; 
  assign auto_sbypass_node_in_in_d_bits_denied = sbypass_auto_node_in_in_d_bits_denied; 
  assign auto_sbypass_node_in_in_d_bits_data = sbypass_auto_node_in_in_d_bits_data; 
  assign auto_sbypass_node_in_in_d_bits_corrupt = sbypass_auto_node_in_in_d_bits_corrupt; 
  assign auto_io_out_c2b_clk = tx_io_c2b_clk; 
  assign auto_io_out_c2b_rst = tx_io_c2b_rst; 
  assign auto_io_out_c2b_send = tx_io_c2b_send; 
  assign auto_io_out_c2b_data = tx_io_c2b_data; 
  assign sbypass_clock = clock; 
  assign sbypass_reset = reset; 
  assign sbypass_auto_node_out_out_a_ready = sinkA_io_a_ready; 
  assign sbypass_auto_node_out_out_d_valid = sourceD_io_d_valid; 
  assign sbypass_auto_node_out_out_d_bits_opcode = sourceD_io_d_bits_opcode; 
  assign sbypass_auto_node_out_out_d_bits_param = sourceD_io_d_bits_param; 
  assign sbypass_auto_node_out_out_d_bits_size = sourceD_io_d_bits_size; 
  assign sbypass_auto_node_out_out_d_bits_source = sourceD_io_d_bits_source; 
  assign sbypass_auto_node_out_out_d_bits_sink = sourceD_io_d_bits_sink; 
  assign sbypass_auto_node_out_out_d_bits_denied = sourceD_io_d_bits_denied; 
  assign sbypass_auto_node_out_out_d_bits_data = sourceD_io_d_bits_data; 
  assign sbypass_auto_node_out_out_d_bits_corrupt = sourceD_io_d_bits_corrupt; 
  assign sbypass_auto_node_in_in_a_valid = auto_sbypass_node_in_in_a_valid; 
  assign sbypass_auto_node_in_in_a_bits_opcode = auto_sbypass_node_in_in_a_bits_opcode; 
  assign sbypass_auto_node_in_in_a_bits_param = auto_sbypass_node_in_in_a_bits_param; 
  assign sbypass_auto_node_in_in_a_bits_size = auto_sbypass_node_in_in_a_bits_size; 
  assign sbypass_auto_node_in_in_a_bits_source = auto_sbypass_node_in_in_a_bits_source; 
  assign sbypass_auto_node_in_in_a_bits_address = auto_sbypass_node_in_in_a_bits_address; 
  assign sbypass_auto_node_in_in_a_bits_mask = auto_sbypass_node_in_in_a_bits_mask; 
  assign sbypass_auto_node_in_in_a_bits_data = auto_sbypass_node_in_in_a_bits_data; 
  assign sbypass_auto_node_in_in_a_bits_corrupt = auto_sbypass_node_in_in_a_bits_corrupt; 
  assign sbypass_auto_node_in_in_d_ready = auto_sbypass_node_in_in_d_ready; 
  assign sbypass_io_bypass = ResetCatchAndSync_d3_io_sync_reset | ResetCatchAndSync_d3_1_io_sync_reset; 
  assign mbypass_clock = clock; 
  assign mbypass_reset = reset; 
  assign mbypass_auto_in_1_a_valid = sourceA_io_a_valid; 
  assign mbypass_auto_in_1_a_bits_opcode = sourceA_io_a_bits_opcode; 
  assign mbypass_auto_in_1_a_bits_param = sourceA_io_a_bits_param; 
  assign mbypass_auto_in_1_a_bits_size = sourceA_io_a_bits_size; 
  assign mbypass_auto_in_1_a_bits_source = sourceA_io_a_bits_source; 
  assign mbypass_auto_in_1_a_bits_address = sourceA_io_a_bits_address; 
  assign mbypass_auto_in_1_a_bits_mask = sourceA_io_a_bits_mask; 
  assign mbypass_auto_in_1_a_bits_data = sourceA_io_a_bits_data; 
  assign mbypass_auto_in_1_c_valid = sourceC_io_c_valid; 
  assign mbypass_auto_in_1_c_bits_opcode = sourceC_io_c_bits_opcode; 
  assign mbypass_auto_in_1_c_bits_param = sourceC_io_c_bits_param; 
  assign mbypass_auto_in_1_c_bits_size = sourceC_io_c_bits_size; 
  assign mbypass_auto_in_1_c_bits_source = sourceC_io_c_bits_source; 
  assign mbypass_auto_in_1_c_bits_address = sourceC_io_c_bits_address; 
  assign mbypass_auto_in_1_d_ready = sinkD_io_d_ready; 
  assign mbypass_auto_in_1_e_valid = sourceE_io_e_valid; 
  assign mbypass_auto_in_1_e_bits_sink = sourceE_io_e_bits_sink; 
  assign mbypass_auto_in_0_c_valid = buffer_auto_out_c_valid; 
  assign mbypass_auto_in_0_c_bits_opcode = buffer_auto_out_c_bits_opcode; 
  assign mbypass_auto_in_0_c_bits_param = buffer_auto_out_c_bits_param; 
  assign mbypass_auto_in_0_c_bits_size = buffer_auto_out_c_bits_size; 
  assign mbypass_auto_in_0_c_bits_source = buffer_auto_out_c_bits_source; 
  assign mbypass_auto_in_0_c_bits_address = buffer_auto_out_c_bits_address; 
  assign mbypass_auto_in_0_c_bits_corrupt = buffer_auto_out_c_bits_corrupt; 
  assign mbypass_auto_out_a_ready = auto_mbypass_out_a_ready; 
  assign mbypass_auto_out_c_ready = auto_mbypass_out_c_ready; 
  assign mbypass_auto_out_d_valid = auto_mbypass_out_d_valid; 
  assign mbypass_auto_out_d_bits_opcode = auto_mbypass_out_d_bits_opcode; 
  assign mbypass_auto_out_d_bits_param = auto_mbypass_out_d_bits_param; 
  assign mbypass_auto_out_d_bits_size = auto_mbypass_out_d_bits_size; 
  assign mbypass_auto_out_d_bits_source = auto_mbypass_out_d_bits_source; 
  assign mbypass_auto_out_d_bits_sink = auto_mbypass_out_d_bits_sink; 
  assign mbypass_auto_out_d_bits_denied = auto_mbypass_out_d_bits_denied; 
  assign mbypass_auto_out_d_bits_data = auto_mbypass_out_d_bits_data; 
  assign mbypass_auto_out_d_bits_corrupt = auto_mbypass_out_d_bits_corrupt; 
  assign mbypass_auto_out_e_ready = auto_mbypass_out_e_ready; 
  assign mbypass_io_bypass = ResetCatchAndSync_d3_io_sync_reset | ResetCatchAndSync_d3_1_io_sync_reset; 
  assign buffer_clock = clock; 
  assign buffer_reset = reset; 
  assign buffer_auto_out_c_ready = mbypass_auto_in_0_c_ready; 
  assign buffer_auto_out_d_valid = mbypass_auto_in_0_d_valid; 
  assign buffer_auto_out_d_bits_opcode = mbypass_auto_in_0_d_bits_opcode; 
  assign buffer_auto_out_d_bits_param = mbypass_auto_in_0_d_bits_param; 
  assign buffer_auto_out_d_bits_size = mbypass_auto_in_0_d_bits_size; 
  assign buffer_auto_out_d_bits_source = mbypass_auto_in_0_d_bits_source; 
  assign buffer_auto_out_d_bits_sink = mbypass_auto_in_0_d_bits_sink; 
  assign buffer_auto_out_d_bits_denied = mbypass_auto_in_0_d_bits_denied; 
  assign buffer_auto_out_d_bits_corrupt = mbypass_auto_in_0_d_bits_corrupt; 
  assign TLMonitor_clock = clock; 
  assign TLMonitor_reset = reset; 
  assign TLMonitor_io_in_a_ready = sinkA_io_a_ready; 
  assign TLMonitor_io_in_a_valid = sbypass_auto_node_out_out_a_valid; 
  assign TLMonitor_io_in_a_bits_opcode = sbypass_auto_node_out_out_a_bits_opcode; 
  assign TLMonitor_io_in_a_bits_param = sbypass_auto_node_out_out_a_bits_param; 
  assign TLMonitor_io_in_a_bits_size = sbypass_auto_node_out_out_a_bits_size; 
  assign TLMonitor_io_in_a_bits_source = sbypass_auto_node_out_out_a_bits_source; 
  assign TLMonitor_io_in_a_bits_address = sbypass_auto_node_out_out_a_bits_address; 
  assign TLMonitor_io_in_a_bits_mask = sbypass_auto_node_out_out_a_bits_mask; 
  assign TLMonitor_io_in_a_bits_corrupt = sbypass_auto_node_out_out_a_bits_corrupt; 
  assign TLMonitor_io_in_bvalid = sourceB_io_bvalid; 
  assign TLMonitor_io_in_d_ready = sbypass_auto_node_out_out_d_ready; 
  assign TLMonitor_io_in_d_valid = sourceD_io_d_valid; 
  assign TLMonitor_io_in_d_bits_opcode = sourceD_io_d_bits_opcode; 
  assign TLMonitor_io_in_d_bits_param = sourceD_io_d_bits_param; 
  assign TLMonitor_io_in_d_bits_size = sourceD_io_d_bits_size; 
  assign TLMonitor_io_in_d_bits_source = sourceD_io_d_bits_source; 
  assign TLMonitor_io_in_d_bits_sink = sourceD_io_d_bits_sink; 
  assign TLMonitor_io_in_d_bits_denied = sourceD_io_d_bits_denied; 
  assign TLMonitor_io_in_d_bits_corrupt = sourceD_io_d_bits_corrupt; 
  assign sinkA_clock = clock; 
  assign sinkA_reset = reset; 
  assign sinkA_io_a_valid = sbypass_auto_node_out_out_a_valid; 
  assign sinkA_io_a_bits_opcode = sbypass_auto_node_out_out_a_bits_opcode; 
  assign sinkA_io_a_bits_param = sbypass_auto_node_out_out_a_bits_param; 
  assign sinkA_io_a_bits_size = sbypass_auto_node_out_out_a_bits_size; 
  assign sinkA_io_a_bits_source = sbypass_auto_node_out_out_a_bits_source; 
  assign sinkA_io_a_bits_address = sbypass_auto_node_out_out_a_bits_address; 
  assign sinkA_io_a_bits_mask = sbypass_auto_node_out_out_a_bits_mask; 
  assign sinkA_io_a_bits_data = sbypass_auto_node_out_out_a_bits_data; 
  assign sinkA_io_q_ready = tx_io_sa_ready; 
  assign sinkB_clock = clock; 
  assign sinkB_reset = reset; 
  assign sinkB_io_q_ready = tx_io_sb_ready; 
  assign sinkC_clock = clock; 
  assign sinkC_reset = reset; 
  assign sinkC_io_q_ready = tx_io_sc_ready; 
  assign sinkD_clock = clock; 
  assign sinkD_reset = reset; 
  assign sinkD_io_d_valid = mbypass_auto_in_1_d_valid; 
  assign sinkD_io_d_bits_opcode = mbypass_auto_in_1_d_bits_opcode; 
  assign sinkD_io_d_bits_param = mbypass_auto_in_1_d_bits_param; 
  assign sinkD_io_d_bits_size = mbypass_auto_in_1_d_bits_size; 
  assign sinkD_io_d_bits_source = mbypass_auto_in_1_d_bits_source; 
  assign sinkD_io_d_bits_sink = mbypass_auto_in_1_d_bits_sink; 
  assign sinkD_io_d_bits_denied = mbypass_auto_in_1_d_bits_denied; 
  assign sinkD_io_d_bits_data = mbypass_auto_in_1_d_bits_data; 
  assign sinkD_io_q_ready = tx_io_sd_ready; 
  assign sinkD_io_a_clSource = sourceA_io_d_clSource; 
  assign sinkD_io_c_clSource = sourceC_io_d_clSource; 
  assign sinkE_io_d_clSink = sourceD_io_e_clSink; 
  assign sourceA_clock = clock; 
  assign sourceA_reset = reset; 
  assign sourceA_io_a_ready = mbypass_auto_in_1_a_ready; 
  assign sourceA_io_q_valid = AsyncQueueSink_io_deq_valid; 
  assign sourceA_io_q_bits = AsyncQueueSink_io_deq_bits; 
  assign sourceA_io_d_tlSource_valid = sinkD_io_a_tlSource_valid; 
  assign sourceA_io_d_tlSource_bits = sinkD_io_a_tlSource_bits; 
  assign sourceB_clock = clock; 
  assign sourceB_reset = reset; 
  assign sourceB_io_q_valid = AsyncQueueSink_1_io_deq_valid; 
  assign sourceB_io_q_bits = AsyncQueueSink_1_io_deq_bits; 
  assign sourceC_clock = clock; 
  assign sourceC_reset = reset; 
  assign sourceC_io_c_ready = mbypass_auto_in_1_c_ready; 
  assign sourceC_io_q_valid = AsyncQueueSink_2_io_deq_valid; 
  assign sourceC_io_q_bits = AsyncQueueSink_2_io_deq_bits; 
  assign sourceC_io_d_tlSource_valid = sinkD_io_c_tlSource_valid; 
  assign sourceC_io_d_tlSource_bits = sinkD_io_c_tlSource_bits; 
  assign sourceD_clock = clock; 
  assign sourceD_reset = reset; 
  assign sourceD_io_d_ready = sbypass_auto_node_out_out_d_ready; 
  assign sourceD_io_q_valid = AsyncQueueSink_3_io_deq_valid; 
  assign sourceD_io_q_bits = AsyncQueueSink_3_io_deq_bits; 
  assign sourceE_io_e_ready = mbypass_auto_in_1_e_ready; 
  assign sourceE_io_q_valid = AsyncQueueSink_4_io_deq_valid; 
  assign sourceE_io_q_bits = AsyncQueueSink_4_io_deq_bits; 
  assign rx_clock = auto_io_out_b2c_clk; 
  assign rx_reset = AsyncResetReg_q; 
  assign rx_io_b2c_send = auto_io_out_b2c_send; 
  assign rx_io_b2c_data = auto_io_out_b2c_data; 
  assign rx_io_a_ridx = AsyncQueueSink_io_async_ridx; 
  assign rx_io_a_safe_ridx_valid = AsyncQueueSink_io_async_safe_ridx_valid; 
  assign rx_io_a_safe_sink_reset_n = AsyncQueueSink_io_async_safe_sink_reset_n; 
  assign rx_io_bridx = AsyncQueueSink_1_io_async_ridx; 
  assign rx_io_bsafe_ridx_valid = AsyncQueueSink_1_io_async_safe_ridx_valid; 
  assign rx_io_bsafe_sink_reset_n = AsyncQueueSink_1_io_async_safe_sink_reset_n; 
  assign rx_io_c_ridx = AsyncQueueSink_2_io_async_ridx; 
  assign rx_io_c_safe_ridx_valid = AsyncQueueSink_2_io_async_safe_ridx_valid; 
  assign rx_io_c_safe_sink_reset_n = AsyncQueueSink_2_io_async_safe_sink_reset_n; 
  assign rx_io_d_ridx = AsyncQueueSink_3_io_async_ridx; 
  assign rx_io_d_safe_ridx_valid = AsyncQueueSink_3_io_async_safe_ridx_valid; 
  assign rx_io_d_safe_sink_reset_n = AsyncQueueSink_3_io_async_safe_sink_reset_n; 
  assign rx_io_e_ridx = AsyncQueueSink_4_io_async_ridx; 
  assign rx_io_e_safe_ridx_valid = AsyncQueueSink_4_io_async_safe_ridx_valid; 
  assign rx_io_e_safe_sink_reset_n = AsyncQueueSink_4_io_async_safe_sink_reset_n; 
  assign rx_io_rxc_ridx = tx_io_rxc_ridx; 
  assign rx_io_rxc_safe_ridx_valid = tx_io_rxc_safe_ridx_valid; 
  assign rx_io_rxc_safe_sink_reset_n = tx_io_rxc_safe_sink_reset_n; 
  assign rx_io_txc_ridx = tx_io_txc_ridx; 
  assign rx_io_txc_safe_ridx_valid = tx_io_txc_safe_ridx_valid; 
  assign rx_io_txc_safe_sink_reset_n = tx_io_txc_safe_sink_reset_n; 
  assign AsyncResetReg_d = 1'h0; 
  assign AsyncResetReg_en = 1'h1; 
  assign AsyncResetReg_clk = auto_io_out_b2c_clk; 
  assign AsyncResetReg_rst = auto_io_out_b2c_rst; 
  assign AsyncQueueSink_clock = clock; 
  assign AsyncQueueSink_reset = reset; 
  assign AsyncQueueSink_io_deq_ready = sourceA_io_q_ready; 
  assign AsyncQueueSink_io_async_mem_0 = rx_io_a_mem_0; 
  assign AsyncQueueSink_io_async_mem_1 = rx_io_a_mem_1; 
  assign AsyncQueueSink_io_async_mem_2 = rx_io_a_mem_2; 
  assign AsyncQueueSink_io_async_mem_3 = rx_io_a_mem_3; 
  assign AsyncQueueSink_io_async_mem_4 = rx_io_a_mem_4; 
  assign AsyncQueueSink_io_async_mem_5 = rx_io_a_mem_5; 
  assign AsyncQueueSink_io_async_mem_6 = rx_io_a_mem_6; 
  assign AsyncQueueSink_io_async_mem_7 = rx_io_a_mem_7; 
  assign AsyncQueueSink_io_async_widx = rx_io_a_widx; 
  assign AsyncQueueSink_io_async_safe_widx_valid = rx_io_a_safe_widx_valid; 
  assign AsyncQueueSink_io_async_safe_source_reset_n = rx_io_a_safe_source_reset_n; 
  assign AsyncQueueSink_1_clock = clock; 
  assign AsyncQueueSink_1_reset = reset; 
  assign AsyncQueueSink_1_io_deq_ready = 1'h1; 
  assign AsyncQueueSink_1_io_async_mem_0 = rx_io_bmem_0; 
  assign AsyncQueueSink_1_io_async_mem_1 = rx_io_bmem_1; 
  assign AsyncQueueSink_1_io_async_mem_2 = rx_io_bmem_2; 
  assign AsyncQueueSink_1_io_async_mem_3 = rx_io_bmem_3; 
  assign AsyncQueueSink_1_io_async_mem_4 = rx_io_bmem_4; 
  assign AsyncQueueSink_1_io_async_mem_5 = rx_io_bmem_5; 
  assign AsyncQueueSink_1_io_async_mem_6 = rx_io_bmem_6; 
  assign AsyncQueueSink_1_io_async_mem_7 = rx_io_bmem_7; 
  assign AsyncQueueSink_1_io_async_widx = rx_io_bwidx; 
  assign AsyncQueueSink_1_io_async_safe_widx_valid = rx_io_bsafe_widx_valid; 
  assign AsyncQueueSink_1_io_async_safe_source_reset_n = rx_io_bsafe_source_reset_n; 
  assign AsyncQueueSink_2_clock = clock; 
  assign AsyncQueueSink_2_reset = reset; 
  assign AsyncQueueSink_2_io_deq_ready = sourceC_io_q_ready; 
  assign AsyncQueueSink_2_io_async_mem_0 = rx_io_c_mem_0; 
  assign AsyncQueueSink_2_io_async_mem_1 = rx_io_c_mem_1; 
  assign AsyncQueueSink_2_io_async_mem_2 = rx_io_c_mem_2; 
  assign AsyncQueueSink_2_io_async_mem_3 = rx_io_c_mem_3; 
  assign AsyncQueueSink_2_io_async_mem_4 = rx_io_c_mem_4; 
  assign AsyncQueueSink_2_io_async_mem_5 = rx_io_c_mem_5; 
  assign AsyncQueueSink_2_io_async_mem_6 = rx_io_c_mem_6; 
  assign AsyncQueueSink_2_io_async_mem_7 = rx_io_c_mem_7; 
  assign AsyncQueueSink_2_io_async_widx = rx_io_c_widx; 
  assign AsyncQueueSink_2_io_async_safe_widx_valid = rx_io_c_safe_widx_valid; 
  assign AsyncQueueSink_2_io_async_safe_source_reset_n = rx_io_c_safe_source_reset_n; 
  assign AsyncQueueSink_3_clock = clock; 
  assign AsyncQueueSink_3_reset = reset; 
  assign AsyncQueueSink_3_io_deq_ready = sourceD_io_q_ready; 
  assign AsyncQueueSink_3_io_async_mem_0 = rx_io_d_mem_0; 
  assign AsyncQueueSink_3_io_async_mem_1 = rx_io_d_mem_1; 
  assign AsyncQueueSink_3_io_async_mem_2 = rx_io_d_mem_2; 
  assign AsyncQueueSink_3_io_async_mem_3 = rx_io_d_mem_3; 
  assign AsyncQueueSink_3_io_async_mem_4 = rx_io_d_mem_4; 
  assign AsyncQueueSink_3_io_async_mem_5 = rx_io_d_mem_5; 
  assign AsyncQueueSink_3_io_async_mem_6 = rx_io_d_mem_6; 
  assign AsyncQueueSink_3_io_async_mem_7 = rx_io_d_mem_7; 
  assign AsyncQueueSink_3_io_async_widx = rx_io_d_widx; 
  assign AsyncQueueSink_3_io_async_safe_widx_valid = rx_io_d_safe_widx_valid; 
  assign AsyncQueueSink_3_io_async_safe_source_reset_n = rx_io_d_safe_source_reset_n; 
  assign AsyncQueueSink_4_clock = clock; 
  assign AsyncQueueSink_4_reset = reset; 
  assign AsyncQueueSink_4_io_deq_ready = sourceE_io_q_ready; 
  assign AsyncQueueSink_4_io_async_mem_0 = rx_io_e_mem_0; 
  assign AsyncQueueSink_4_io_async_mem_1 = rx_io_e_mem_1; 
  assign AsyncQueueSink_4_io_async_mem_2 = rx_io_e_mem_2; 
  assign AsyncQueueSink_4_io_async_mem_3 = rx_io_e_mem_3; 
  assign AsyncQueueSink_4_io_async_mem_4 = rx_io_e_mem_4; 
  assign AsyncQueueSink_4_io_async_mem_5 = rx_io_e_mem_5; 
  assign AsyncQueueSink_4_io_async_mem_6 = rx_io_e_mem_6; 
  assign AsyncQueueSink_4_io_async_mem_7 = rx_io_e_mem_7; 
  assign AsyncQueueSink_4_io_async_widx = rx_io_e_widx; 
  assign AsyncQueueSink_4_io_async_safe_widx_valid = rx_io_e_safe_widx_valid; 
  assign AsyncQueueSink_4_io_async_safe_source_reset_n = rx_io_e_safe_source_reset_n; 
  assign tx_clock = clock; 
  assign tx_reset = reset; 
  assign tx_io_sa_valid = sinkA_io_q_valid; 
  assign tx_io_sa_bits_data = sinkA_io_q_bits_data; 
  assign tx_io_sa_bits_last = sinkA_io_q_bits_last; 
  assign tx_io_sa_bits_beats = sinkA_io_q_bits_beats; 
  assign tx_io_sb_bits_data = sinkB_io_q_bits_data; 
  assign tx_io_sb_bits_last = sinkB_io_q_bits_last; 
  assign tx_io_sc_bits_data = sinkC_io_q_bits_data; 
  assign tx_io_sc_bits_last = sinkC_io_q_bits_last; 
  assign tx_io_sd_valid = sinkD_io_q_valid; 
  assign tx_io_sd_bits_data = sinkD_io_q_bits_data; 
  assign tx_io_sd_bits_last = sinkD_io_q_bits_last; 
  assign tx_io_sd_bits_beats = sinkD_io_q_bits_beats; 
  assign tx_io_se_bits_data = sinkE_io_q_bits_data; 
  assign tx_io_rxc_mem_0_a = rx_io_rxc_mem_0_a; 
  assign tx_io_rxc_mem_0_b = rx_io_rxc_mem_0_b; 
  assign tx_io_rxc_mem_0_c = rx_io_rxc_mem_0_c; 
  assign tx_io_rxc_mem_0_d = rx_io_rxc_mem_0_d; 
  assign tx_io_rxc_mem_0_e = rx_io_rxc_mem_0_e; 
  assign tx_io_rxc_widx = rx_io_rxc_widx; 
  assign tx_io_rxc_safe_widx_valid = rx_io_rxc_safe_widx_valid; 
  assign tx_io_rxc_safe_source_reset_n = rx_io_rxc_safe_source_reset_n; 
  assign tx_io_txc_mem_0_a = rx_io_txc_mem_0_a; 
  assign tx_io_txc_mem_0_b = rx_io_txc_mem_0_b; 
  assign tx_io_txc_mem_0_c = rx_io_txc_mem_0_c; 
  assign tx_io_txc_mem_0_d = rx_io_txc_mem_0_d; 
  assign tx_io_txc_mem_0_e = rx_io_txc_mem_0_e; 
  assign tx_io_txc_widx = rx_io_txc_widx; 
  assign tx_io_txc_safe_widx_valid = rx_io_txc_safe_widx_valid; 
  assign tx_io_txc_safe_source_reset_n = rx_io_txc_safe_source_reset_n; 
  assign ResetCatchAndSync_d3_clock = clock; 
  assign ResetCatchAndSync_d3_reset = rx_reset; 
  assign ResetCatchAndSync_d3_1_clock = clock; 
  assign ResetCatchAndSync_d3_1_reset = tx_reset; 
endmodule
module dual_HellaFlowQueue( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [31:0] io_enq_bits, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [31:0] io_deq_bits 
);
  wire [10:0] ram_R0_addr; 
  wire  ram_R0_en; 
  wire  ram_R0_clk; 
  wire [31:0] ram_R0_data; 
  wire [10:0] ram_W0_addr; 
  wire  ram_W0_en; 
  wire  ram_W0_clk; 
  wire [31:0] ram_W0_data; 
  wire  _T; 
  reg [10:0] value; 
  reg [31:0] _RAND_0;
  reg [10:0] value_1; 
  reg [31:0] _RAND_1;
  wire  ptr_match; 
  reg  maybe_full; 
  reg [31:0] _RAND_2;
  wire  _T_12; 
  wire  empty; 
  wire  do_flow; 
  wire  _T_1; 
  wire  do_enq; 
  wire  _T_2; 
  wire  do_deq; 
  wire [10:0] _T_6; 
  wire  _T_8; 
  wire [10:0] _T_10; 
  wire  deq_done; 
  wire  _T_11; 
  wire  full; 
  wire [10:0] _T_14; 
  wire  _T_15; 
  wire  atLeastTwo; 
  wire  _T_18; 
  wire  _T_19; 
  wire  _T_20; 
  wire  _T_21; 
  wire [10:0] _T_24; 
  reg  ram_out_valid; 
  reg [31:0] _RAND_3;
  dual_ram ram ( 
    .R0_addr(ram_R0_addr),
    .R0_en(ram_R0_en),
    .R0_clk(ram_R0_clk),
    .R0_data(ram_R0_data),
    .W0_addr(ram_W0_addr),
    .W0_en(ram_W0_en),
    .W0_clk(ram_W0_clk),
    .W0_data(ram_W0_data)
  );
  assign _T = io_enq_ready & io_enq_valid; 
  assign ptr_match = value == value_1; 
  assign _T_12 = maybe_full == 1'h0; 
  assign empty = ptr_match & _T_12; 
  assign do_flow = empty & io_deq_ready; 
  assign _T_1 = do_flow == 1'h0; 
  assign do_enq = _T & _T_1; 
  assign _T_2 = io_deq_ready & io_deq_valid; 
  assign do_deq = _T_2 & _T_1; 
  assign _T_6 = value + 11'h1; 
  assign _T_8 = value_1 == 11'h7ff; 
  assign _T_10 = value_1 + 11'h1; 
  assign deq_done = do_deq & _T_8; 
  assign _T_11 = do_enq != do_deq; 
  assign full = ptr_match & maybe_full; 
  assign _T_14 = value - value_1; 
  assign _T_15 = _T_14 >= 11'h2; 
  assign atLeastTwo = full | _T_15; 
  assign _T_18 = io_deq_valid == 1'h0; 
  assign _T_19 = empty == 1'h0; 
  assign _T_20 = _T_18 & _T_19; 
  assign _T_21 = atLeastTwo | _T_20; 
  assign _T_24 = deq_done ? 11'h0 : _T_10; 
  assign io_enq_ready = full == 1'h0; 
  assign io_deq_valid = empty ? io_enq_valid : ram_out_valid; 
  assign io_deq_bits = empty ? io_enq_bits : ram_R0_data; 
  assign ram_R0_addr = io_deq_valid ? _T_24 : value_1; 
  assign ram_R0_en = io_deq_ready & _T_21; 
  assign ram_R0_clk = clock; 
  assign ram_W0_addr = value; 
  assign ram_W0_en = _T & _T_1; 
  assign ram_W0_clk = clock; 
  assign ram_W0_data = io_enq_bits; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value_1 = _RAND_1[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ram_out_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 11'h0;
    end else begin
      if (do_enq) begin
        value <= _T_6;
      end
    end
    if (reset) begin
      value_1 <= 11'h0;
    end else begin
      if (do_deq) begin
        value_1 <= _T_10;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_11) begin
        maybe_full <= do_enq;
      end
    end
    ram_out_valid <= io_deq_ready & _T_21;
  end
endmodule
module dual_HellaQueue( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [31:0] io_enq_bits, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [31:0] io_deq_bits 
);
  wire  fq_clock; 
  wire  fq_reset; 
  wire  fq_io_enq_ready; 
  wire  fq_io_enq_valid; 
  wire [31:0] fq_io_enq_bits; 
  wire  fq_io_deq_ready; 
  wire  fq_io_deq_valid; 
  wire [31:0] fq_io_deq_bits; 
  wire  Queue_clock; 
  wire  Queue_reset; 
  wire  Queue_io_enq_ready; 
  wire  Queue_io_enq_valid; 
  wire [31:0] Queue_io_enq_bits; 
  wire  Queue_io_deq_ready; 
  wire  Queue_io_deq_valid; 
  wire [31:0] Queue_io_deq_bits; 
  dual_HellaFlowQueue fq ( 
    .clock(fq_clock),
    .reset(fq_reset),
    .io_enq_ready(fq_io_enq_ready),
    .io_enq_valid(fq_io_enq_valid),
    .io_enq_bits(fq_io_enq_bits),
    .io_deq_ready(fq_io_deq_ready),
    .io_deq_valid(fq_io_deq_valid),
    .io_deq_bits(fq_io_deq_bits)
  );
  dual_Queue_9 dual_Queue ( 
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits(Queue_io_enq_bits),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits(Queue_io_deq_bits)
  );
  assign io_enq_ready = fq_io_enq_ready; 
  assign io_deq_valid = Queue_io_deq_valid; 
  assign io_deq_bits = Queue_io_deq_bits; 
  assign fq_clock = clock; 
  assign fq_reset = reset; 
  assign fq_io_enq_valid = io_enq_valid; 
  assign fq_io_enq_bits = io_enq_bits; 
  assign fq_io_deq_ready = Queue_io_enq_ready; 
  assign Queue_clock = clock; 
  assign Queue_reset = reset; 
  assign Queue_io_enq_valid = fq_io_deq_valid; 
  assign Queue_io_enq_bits = fq_io_deq_bits; 
  assign Queue_io_deq_ready = io_deq_ready; 
endmodule
module dual_MasterMux( 
  input         clock, 
  input         reset, 
  output        auto_in_1_a_ready, 
  input         auto_in_1_a_valid, 
  input  [2:0]  auto_in_1_a_bits_opcode, 
  input  [2:0]  auto_in_1_a_bits_param, 
  input  [3:0]  auto_in_1_a_bits_size, 
  input  [5:0]  auto_in_1_a_bits_source, 
  input  [31:0] auto_in_1_a_bits_address, 
  input  [3:0]  auto_in_1_a_bits_mask, 
  input  [31:0] auto_in_1_a_bits_data, 
  output        auto_in_1_c_ready, 
  input         auto_in_1_c_valid, 
  input  [2:0]  auto_in_1_c_bits_opcode, 
  input  [2:0]  auto_in_1_c_bits_param, 
  input  [3:0]  auto_in_1_c_bits_size, 
  input  [5:0]  auto_in_1_c_bits_source, 
  input  [31:0] auto_in_1_c_bits_address, 
  input         auto_in_1_d_ready, 
  output        auto_in_1_d_valid, 
  output [2:0]  auto_in_1_d_bits_opcode, 
  output [1:0]  auto_in_1_d_bits_param, 
  output [3:0]  auto_in_1_d_bits_size, 
  output [5:0]  auto_in_1_d_bits_source, 
  output        auto_in_1_d_bits_sink, 
  output        auto_in_1_d_bits_denied, 
  output [31:0] auto_in_1_d_bits_data, 
  output        auto_in_1_e_ready, 
  input         auto_in_1_e_valid, 
  input         auto_in_1_e_bits_sink, 
  output        auto_in_0_c_ready, 
  input         auto_in_0_c_valid, 
  input  [2:0]  auto_in_0_c_bits_opcode, 
  input  [2:0]  auto_in_0_c_bits_param, 
  input  [3:0]  auto_in_0_c_bits_size, 
  input         auto_in_0_c_bits_source, 
  input  [31:0] auto_in_0_c_bits_address, 
  input         auto_in_0_c_bits_corrupt, 
  output        auto_in_0_d_valid, 
  output [2:0]  auto_in_0_d_bits_opcode, 
  output [1:0]  auto_in_0_d_bits_param, 
  output [3:0]  auto_in_0_d_bits_size, 
  output        auto_in_0_d_bits_source, 
  output        auto_in_0_d_bits_sink, 
  output        auto_in_0_d_bits_denied, 
  output        auto_in_0_d_bits_corrupt, 
  input         auto_out_a_ready, 
  output        auto_out_a_valid, 
  output [2:0]  auto_out_a_bits_opcode, 
  output [2:0]  auto_out_a_bits_param, 
  output [3:0]  auto_out_a_bits_size, 
  output [5:0]  auto_out_a_bits_source, 
  output [31:0] auto_out_a_bits_address, 
  output [3:0]  auto_out_a_bits_mask, 
  output [31:0] auto_out_a_bits_data, 
  input         auto_out_c_ready, 
  output        auto_out_c_valid, 
  output [2:0]  auto_out_c_bits_opcode, 
  output [2:0]  auto_out_c_bits_param, 
  output [3:0]  auto_out_c_bits_size, 
  output [5:0]  auto_out_c_bits_source, 
  output [31:0] auto_out_c_bits_address, 
  output        auto_out_c_bits_corrupt, 
  output        auto_out_d_ready, 
  input         auto_out_d_valid, 
  input  [2:0]  auto_out_d_bits_opcode, 
  input  [1:0]  auto_out_d_bits_param, 
  input  [3:0]  auto_out_d_bits_size, 
  input  [5:0]  auto_out_d_bits_source, 
  input         auto_out_d_bits_sink, 
  input         auto_out_d_bits_denied, 
  input  [31:0] auto_out_d_bits_data, 
  input         auto_out_d_bits_corrupt, 
  input         auto_out_e_ready, 
  output        auto_out_e_valid, 
  output        auto_out_e_bits_sink, 
  input         io_bypass 
);
  wire  TLMonitor_clock; 
  wire  TLMonitor_reset; 
  wire  TLMonitor_io_in_c_ready; 
  wire  TLMonitor_io_in_c_valid; 
  wire [2:0] TLMonitor_io_in_c_bits_opcode; 
  wire [2:0] TLMonitor_io_in_c_bits_param; 
  wire [3:0] TLMonitor_io_in_c_bits_size; 
  wire  TLMonitor_io_in_c_bits_source; 
  wire [31:0] TLMonitor_io_in_c_bits_address; 
  wire  TLMonitor_io_in_c_bits_corrupt; 
  wire  TLMonitor_io_in_d_valid; 
  wire [2:0] TLMonitor_io_in_d_bits_opcode; 
  wire [1:0] TLMonitor_io_in_d_bits_param; 
  wire [3:0] TLMonitor_io_in_d_bits_size; 
  wire  TLMonitor_io_in_d_bits_source; 
  wire  TLMonitor_io_in_d_bits_sink; 
  wire  TLMonitor_io_in_d_bits_denied; 
  wire  TLMonitor_io_in_d_bits_corrupt; 
  wire  TLMonitor_1_clock; 
  wire  TLMonitor_1_reset; 
  wire  TLMonitor_1_io_in_a_ready; 
  wire  TLMonitor_1_io_in_a_valid; 
  wire [2:0] TLMonitor_1_io_in_a_bits_opcode; 
  wire [2:0] TLMonitor_1_io_in_a_bits_param; 
  wire [3:0] TLMonitor_1_io_in_a_bits_size; 
  wire [5:0] TLMonitor_1_io_in_a_bits_source; 
  wire [31:0] TLMonitor_1_io_in_a_bits_address; 
  wire [3:0] TLMonitor_1_io_in_a_bits_mask; 
  wire  TLMonitor_1_io_in_c_ready; 
  wire  TLMonitor_1_io_in_c_valid; 
  wire [2:0] TLMonitor_1_io_in_c_bits_opcode; 
  wire [2:0] TLMonitor_1_io_in_c_bits_param; 
  wire [3:0] TLMonitor_1_io_in_c_bits_size; 
  wire [5:0] TLMonitor_1_io_in_c_bits_source; 
  wire [31:0] TLMonitor_1_io_in_c_bits_address; 
  wire  TLMonitor_1_io_in_d_ready; 
  wire  TLMonitor_1_io_in_d_valid; 
  wire [2:0] TLMonitor_1_io_in_d_bits_opcode; 
  wire [1:0] TLMonitor_1_io_in_d_bits_param; 
  wire [3:0] TLMonitor_1_io_in_d_bits_size; 
  wire [5:0] TLMonitor_1_io_in_d_bits_source; 
  wire  TLMonitor_1_io_in_d_bits_sink; 
  wire  TLMonitor_1_io_in_d_bits_denied; 
  wire  TLMonitor_1_io_in_d_bits_corrupt; 
  wire  TLMonitor_1_io_in_e_ready; 
  wire  TLMonitor_1_io_in_e_valid; 
  wire  TLMonitor_1_io_in_e_bits_sink; 
  reg  bypass; 
  reg [31:0] _RAND_0;
  reg [7:0] flight; 
  reg [31:0] _RAND_1;
  wire  _T_175; 
  reg [5:0] _T_185; 
  reg [31:0] _RAND_2;
  wire  _T_188; 
  wire  stall; 
  wire  _T_203; 
  wire  _T_204; 
  wire  out_a_valid; 
  wire  _T_12; 
  wire [3:0] out_a_bits_size; 
  wire [22:0] _T_14; 
  wire [7:0] _T_15; 
  wire [7:0] _T_16; 
  wire [5:0] _T_17; 
  wire [2:0] out_a_bits_opcode; 
  wire  _T_18; 
  wire  _T_19; 
  reg [5:0] _T_21; 
  reg [31:0] _RAND_3;
  wire [5:0] _T_23; 
  wire  _T_24; 
  wire  out_c_valid; 
  wire  _T_52; 
  wire [3:0] out_c_bits_size; 
  wire [22:0] _T_54; 
  wire [7:0] _T_55; 
  wire [7:0] _T_56; 
  wire [5:0] _T_57; 
  wire [2:0] out_c_bits_opcode; 
  wire  _T_58; 
  wire [5:0] _T_59; 
  reg [5:0] _T_60; 
  reg [31:0] _RAND_4;
  wire [5:0] _T_62; 
  wire  _T_63; 
  wire  _T_64; 
  wire  _T_65; 
  wire  _T_66; 
  wire  out_d_ready; 
  wire  _T_71; 
  wire [22:0] _T_73; 
  wire [7:0] _T_74; 
  wire [7:0] _T_75; 
  wire [5:0] _T_76; 
  wire  _T_77; 
  wire [5:0] _T_78; 
  reg [5:0] _T_79; 
  reg [31:0] _RAND_5;
  wire [5:0] _T_81; 
  wire  _T_82; 
  wire  _T_83; 
  wire  _T_84; 
  wire  _T_85; 
  wire  out_e_valid; 
  wire  _T_90; 
  wire  _T_102; 
  wire  _T_103; 
  wire  _T_104; 
  wire  _T_106; 
  wire  _T_108; 
  wire  _T_109; 
  wire  _T_110; 
  wire  _T_111; 
  wire  _T_112; 
  wire  _T_113; 
  wire  _T_115; 
  wire  _T_121; 
  wire  _T_122; 
  wire  _T_124; 
  wire  _T_125; 
  wire [4:0] _T_132; 
  wire  _T_140; 
  wire  _T_141; 
  wire  _T_143; 
  wire [4:0] _T_151; 
  wire  _T_152; 
  wire  _T_153; 
  wire  _T_154; 
  wire  _T_155; 
  wire  _T_156; 
  wire [1:0] _T_157; 
  wire [1:0] _T_158; 
  wire [1:0] _GEN_7; 
  wire [2:0] _T_159; 
  wire [2:0] _GEN_8; 
  wire [3:0] _T_160; 
  wire [7:0] _GEN_9; 
  wire [7:0] _T_162; 
  wire  _T_163; 
  wire  _T_164; 
  wire  _T_165; 
  wire  _T_166; 
  wire  _T_167; 
  wire [1:0] _T_168; 
  wire [1:0] _T_169; 
  wire [1:0] _GEN_10; 
  wire [2:0] _T_170; 
  wire [2:0] _GEN_11; 
  wire [3:0] _T_171; 
  wire [7:0] _GEN_12; 
  wire [7:0] next_flight; 
  wire  _T_174; 
  wire [5:0] _T_187; 
  wire  _T_197; 
  wire  _T_201; 
  wire [5:0] _T_221_source; 
  dual_TLMonitor_5 dual_TLMonitor ( 
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_c_ready(TLMonitor_io_in_c_ready),
    .io_in_c_valid(TLMonitor_io_in_c_valid),
    .io_in_c_bits_opcode(TLMonitor_io_in_c_bits_opcode),
    .io_in_c_bits_param(TLMonitor_io_in_c_bits_param),
    .io_in_c_bits_size(TLMonitor_io_in_c_bits_size),
    .io_in_c_bits_source(TLMonitor_io_in_c_bits_source),
    .io_in_c_bits_address(TLMonitor_io_in_c_bits_address),
    .io_in_c_bits_corrupt(TLMonitor_io_in_c_bits_corrupt),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt)
  );
  dual_TLMonitor_6 dual_TLMonitor_1 ( 
    .clock(TLMonitor_1_clock),
    .reset(TLMonitor_1_reset),
    .io_in_a_ready(TLMonitor_1_io_in_a_ready),
    .io_in_a_valid(TLMonitor_1_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_1_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_1_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_1_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_1_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_1_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_1_io_in_a_bits_mask),
    .io_in_c_ready(TLMonitor_1_io_in_c_ready),
    .io_in_c_valid(TLMonitor_1_io_in_c_valid),
    .io_in_c_bits_opcode(TLMonitor_1_io_in_c_bits_opcode),
    .io_in_c_bits_param(TLMonitor_1_io_in_c_bits_param),
    .io_in_c_bits_size(TLMonitor_1_io_in_c_bits_size),
    .io_in_c_bits_source(TLMonitor_1_io_in_c_bits_source),
    .io_in_c_bits_address(TLMonitor_1_io_in_c_bits_address),
    .io_in_d_ready(TLMonitor_1_io_in_d_ready),
    .io_in_d_valid(TLMonitor_1_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_1_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_1_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_1_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_1_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_1_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_1_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_1_io_in_d_bits_corrupt),
    .io_in_e_ready(TLMonitor_1_io_in_e_ready),
    .io_in_e_valid(TLMonitor_1_io_in_e_valid),
    .io_in_e_bits_sink(TLMonitor_1_io_in_e_bits_sink)
  );
  assign _T_175 = bypass != io_bypass; 
  assign _T_188 = _T_185 == 6'h0; 
  assign stall = _T_175 & _T_188; 
  assign _T_203 = stall == 1'h0; 
  assign _T_204 = bypass ? 1'h0 : auto_in_1_a_valid; 
  assign out_a_valid = _T_203 & _T_204; 
  assign _T_12 = auto_out_a_ready & out_a_valid; 
  assign out_a_bits_size = bypass ? 4'h0 : auto_in_1_a_bits_size; 
  assign _T_14 = 23'hff << out_a_bits_size; 
  assign _T_15 = _T_14[7:0]; 
  assign _T_16 = ~ _T_15; 
  assign _T_17 = _T_16[7:2]; 
  assign out_a_bits_opcode = bypass ? 3'h0 : auto_in_1_a_bits_opcode; 
  assign _T_18 = out_a_bits_opcode[2]; 
  assign _T_19 = _T_18 == 1'h0; 
  assign _T_23 = _T_21 - 6'h1; 
  assign _T_24 = _T_21 == 6'h0; 
  assign out_c_valid = bypass ? auto_in_0_c_valid : auto_in_1_c_valid; 
  assign _T_52 = auto_out_c_ready & out_c_valid; 
  assign out_c_bits_size = bypass ? auto_in_0_c_bits_size : auto_in_1_c_bits_size; 
  assign _T_54 = 23'hff << out_c_bits_size; 
  assign _T_55 = _T_54[7:0]; 
  assign _T_56 = ~ _T_55; 
  assign _T_57 = _T_56[7:2]; 
  assign out_c_bits_opcode = bypass ? auto_in_0_c_bits_opcode : auto_in_1_c_bits_opcode; 
  assign _T_58 = out_c_bits_opcode[0]; 
  assign _T_59 = _T_58 ? _T_57 : 6'h0; 
  assign _T_62 = _T_60 - 6'h1; 
  assign _T_63 = _T_60 == 6'h0; 
  assign _T_64 = _T_60 == 6'h1; 
  assign _T_65 = _T_59 == 6'h0; 
  assign _T_66 = _T_64 | _T_65; 
  assign out_d_ready = bypass ? 1'h1 : auto_in_1_d_ready; 
  assign _T_71 = out_d_ready & auto_out_d_valid; 
  assign _T_73 = 23'hff << auto_out_d_bits_size; 
  assign _T_74 = _T_73[7:0]; 
  assign _T_75 = ~ _T_74; 
  assign _T_76 = _T_75[7:2]; 
  assign _T_77 = auto_out_d_bits_opcode[0]; 
  assign _T_78 = _T_77 ? _T_76 : 6'h0; 
  assign _T_81 = _T_79 - 6'h1; 
  assign _T_82 = _T_79 == 6'h0; 
  assign _T_83 = _T_79 == 6'h1; 
  assign _T_84 = _T_78 == 6'h0; 
  assign _T_85 = _T_83 | _T_84; 
  assign out_e_valid = bypass ? 1'h0 : auto_in_1_e_valid; 
  assign _T_90 = auto_out_e_ready & out_e_valid; 
  assign _T_102 = out_c_bits_opcode[2]; 
  assign _T_103 = out_c_bits_opcode[1]; 
  assign _T_104 = _T_102 & _T_103; 
  assign _T_106 = _T_102 == 1'h0; 
  assign _T_108 = _T_103 == 1'h0; 
  assign _T_109 = _T_106 | _T_108; 
  assign _T_110 = auto_out_d_bits_opcode[2]; 
  assign _T_111 = auto_out_d_bits_opcode[1]; 
  assign _T_112 = _T_111 == 1'h0; 
  assign _T_113 = _T_110 & _T_112; 
  assign _T_115 = _T_12 & _T_24; 
  assign _T_121 = _T_52 & _T_63; 
  assign _T_122 = _T_121 & _T_104; 
  assign _T_124 = _T_71 & _T_82; 
  assign _T_125 = _T_124 & _T_113; 
  assign _T_132 = {_T_115,_T_125,1'h0,_T_122,1'h0}; 
  assign _T_140 = _T_52 & _T_66; 
  assign _T_141 = _T_140 & _T_109; 
  assign _T_143 = _T_71 & _T_85; 
  assign _T_151 = {1'h0,_T_143,1'h0,_T_141,_T_90}; 
  assign _T_152 = _T_132[0]; 
  assign _T_153 = _T_132[1]; 
  assign _T_154 = _T_132[2]; 
  assign _T_155 = _T_132[3]; 
  assign _T_156 = _T_132[4]; 
  assign _T_157 = _T_152 + _T_153; 
  assign _T_158 = _T_155 + _T_156; 
  assign _GEN_7 = {{1'd0}, _T_154}; 
  assign _T_159 = _GEN_7 + _T_158; 
  assign _GEN_8 = {{1'd0}, _T_157}; 
  assign _T_160 = _GEN_8 + _T_159; 
  assign _GEN_9 = {{4'd0}, _T_160}; 
  assign _T_162 = flight + _GEN_9; 
  assign _T_163 = _T_151[0]; 
  assign _T_164 = _T_151[1]; 
  assign _T_165 = _T_151[2]; 
  assign _T_166 = _T_151[3]; 
  assign _T_167 = _T_151[4]; 
  assign _T_168 = _T_163 + _T_164; 
  assign _T_169 = _T_166 + _T_167; 
  assign _GEN_10 = {{1'd0}, _T_165}; 
  assign _T_170 = _GEN_10 + _T_169; 
  assign _GEN_11 = {{1'd0}, _T_168}; 
  assign _T_171 = _GEN_11 + _T_170; 
  assign _GEN_12 = {{4'd0}, _T_171}; 
  assign next_flight = _T_162 - _GEN_12; 
  assign _T_174 = next_flight == 8'h0; 
  assign _T_187 = _T_185 - 6'h1; 
  assign _T_197 = _T_203 & auto_out_a_ready; 
  assign _T_201 = bypass == 1'h0; 
  assign _T_221_source = {{5'd0}, auto_in_0_c_bits_source}; 
  assign auto_in_1_a_ready = _T_197 & _T_201; 
  assign auto_in_1_c_ready = auto_out_c_ready & _T_201; 
  assign auto_in_1_d_valid = auto_out_d_valid & _T_201; 
  assign auto_in_1_d_bits_opcode = auto_out_d_bits_opcode; 
  assign auto_in_1_d_bits_param = auto_out_d_bits_param; 
  assign auto_in_1_d_bits_size = auto_out_d_bits_size; 
  assign auto_in_1_d_bits_source = auto_out_d_bits_source; 
  assign auto_in_1_d_bits_sink = auto_out_d_bits_sink; 
  assign auto_in_1_d_bits_denied = auto_out_d_bits_denied; 
  assign auto_in_1_d_bits_data = auto_out_d_bits_data; 
  assign auto_in_1_e_ready = auto_out_e_ready & _T_201; 
  assign auto_in_0_c_ready = auto_out_c_ready & bypass; 
  assign auto_in_0_d_valid = auto_out_d_valid & bypass; 
  assign auto_in_0_d_bits_opcode = auto_out_d_bits_opcode; 
  assign auto_in_0_d_bits_param = auto_out_d_bits_param; 
  assign auto_in_0_d_bits_size = auto_out_d_bits_size; 
  assign auto_in_0_d_bits_source = auto_out_d_bits_source[0]; 
  assign auto_in_0_d_bits_sink = auto_out_d_bits_sink; 
  assign auto_in_0_d_bits_denied = auto_out_d_bits_denied; 
  assign auto_in_0_d_bits_corrupt = auto_out_d_bits_corrupt; 
  assign auto_out_a_valid = _T_203 & _T_204; 
  assign auto_out_a_bits_opcode = bypass ? 3'h0 : auto_in_1_a_bits_opcode; 
  assign auto_out_a_bits_param = bypass ? 3'h0 : auto_in_1_a_bits_param; 
  assign auto_out_a_bits_size = bypass ? 4'h0 : auto_in_1_a_bits_size; 
  assign auto_out_a_bits_source = bypass ? 6'h0 : auto_in_1_a_bits_source; 
  assign auto_out_a_bits_address = bypass ? 32'h0 : auto_in_1_a_bits_address; 
  assign auto_out_a_bits_mask = bypass ? 4'h0 : auto_in_1_a_bits_mask; 
  assign auto_out_a_bits_data = bypass ? 32'h0 : auto_in_1_a_bits_data; 
  assign auto_out_c_valid = bypass ? auto_in_0_c_valid : auto_in_1_c_valid; 
  assign auto_out_c_bits_opcode = bypass ? auto_in_0_c_bits_opcode : auto_in_1_c_bits_opcode; 
  assign auto_out_c_bits_param = bypass ? auto_in_0_c_bits_param : auto_in_1_c_bits_param; 
  assign auto_out_c_bits_size = bypass ? auto_in_0_c_bits_size : auto_in_1_c_bits_size; 
  assign auto_out_c_bits_source = bypass ? _T_221_source : auto_in_1_c_bits_source; 
  assign auto_out_c_bits_address = bypass ? auto_in_0_c_bits_address : auto_in_1_c_bits_address; 
  assign auto_out_c_bits_corrupt = bypass ? auto_in_0_c_bits_corrupt : 1'h0; 
  assign auto_out_d_ready = bypass ? 1'h1 : auto_in_1_d_ready; 
  assign auto_out_e_valid = bypass ? 1'h0 : auto_in_1_e_valid; 
  assign auto_out_e_bits_sink = bypass ? 1'h0 : auto_in_1_e_bits_sink; 
  assign TLMonitor_clock = clock; 
  assign TLMonitor_reset = reset; 
  assign TLMonitor_io_in_c_ready = auto_out_c_ready & bypass; 
  assign TLMonitor_io_in_c_valid = auto_in_0_c_valid; 
  assign TLMonitor_io_in_c_bits_opcode = auto_in_0_c_bits_opcode; 
  assign TLMonitor_io_in_c_bits_param = auto_in_0_c_bits_param; 
  assign TLMonitor_io_in_c_bits_size = auto_in_0_c_bits_size; 
  assign TLMonitor_io_in_c_bits_source = auto_in_0_c_bits_source; 
  assign TLMonitor_io_in_c_bits_address = auto_in_0_c_bits_address; 
  assign TLMonitor_io_in_c_bits_corrupt = auto_in_0_c_bits_corrupt; 
  assign TLMonitor_io_in_d_valid = auto_out_d_valid & bypass; 
  assign TLMonitor_io_in_d_bits_opcode = auto_out_d_bits_opcode; 
  assign TLMonitor_io_in_d_bits_param = auto_out_d_bits_param; 
  assign TLMonitor_io_in_d_bits_size = auto_out_d_bits_size; 
  assign TLMonitor_io_in_d_bits_source = auto_out_d_bits_source[0]; 
  assign TLMonitor_io_in_d_bits_sink = auto_out_d_bits_sink; 
  assign TLMonitor_io_in_d_bits_denied = auto_out_d_bits_denied; 
  assign TLMonitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; 
  assign TLMonitor_1_clock = clock; 
  assign TLMonitor_1_reset = reset; 
  assign TLMonitor_1_io_in_a_ready = _T_197 & _T_201; 
  assign TLMonitor_1_io_in_a_valid = auto_in_1_a_valid; 
  assign TLMonitor_1_io_in_a_bits_opcode = auto_in_1_a_bits_opcode; 
  assign TLMonitor_1_io_in_a_bits_param = auto_in_1_a_bits_param; 
  assign TLMonitor_1_io_in_a_bits_size = auto_in_1_a_bits_size; 
  assign TLMonitor_1_io_in_a_bits_source = auto_in_1_a_bits_source; 
  assign TLMonitor_1_io_in_a_bits_address = auto_in_1_a_bits_address; 
  assign TLMonitor_1_io_in_a_bits_mask = auto_in_1_a_bits_mask; 
  assign TLMonitor_1_io_in_c_ready = auto_out_c_ready & _T_201; 
  assign TLMonitor_1_io_in_c_valid = auto_in_1_c_valid; 
  assign TLMonitor_1_io_in_c_bits_opcode = auto_in_1_c_bits_opcode; 
  assign TLMonitor_1_io_in_c_bits_param = auto_in_1_c_bits_param; 
  assign TLMonitor_1_io_in_c_bits_size = auto_in_1_c_bits_size; 
  assign TLMonitor_1_io_in_c_bits_source = auto_in_1_c_bits_source; 
  assign TLMonitor_1_io_in_c_bits_address = auto_in_1_c_bits_address; 
  assign TLMonitor_1_io_in_d_ready = auto_in_1_d_ready; 
  assign TLMonitor_1_io_in_d_valid = auto_out_d_valid & _T_201; 
  assign TLMonitor_1_io_in_d_bits_opcode = auto_out_d_bits_opcode; 
  assign TLMonitor_1_io_in_d_bits_param = auto_out_d_bits_param; 
  assign TLMonitor_1_io_in_d_bits_size = auto_out_d_bits_size; 
  assign TLMonitor_1_io_in_d_bits_source = auto_out_d_bits_source; 
  assign TLMonitor_1_io_in_d_bits_sink = auto_out_d_bits_sink; 
  assign TLMonitor_1_io_in_d_bits_denied = auto_out_d_bits_denied; 
  assign TLMonitor_1_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; 
  assign TLMonitor_1_io_in_e_ready = auto_out_e_ready & _T_201; 
  assign TLMonitor_1_io_in_e_valid = auto_in_1_e_valid; 
  assign TLMonitor_1_io_in_e_bits_sink = auto_in_1_e_bits_sink; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bypass = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  flight = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_185 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_21 = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_60 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_79 = _RAND_5[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      bypass <= io_bypass;
    end else begin
      if (_T_174) begin
        bypass <= io_bypass;
      end
    end
    if (reset) begin
      flight <= 8'h0;
    end else begin
      flight <= next_flight;
    end
    if (reset) begin
      _T_185 <= 6'h0;
    end else begin
      if (_T_12) begin
        if (_T_188) begin
          if (_T_19) begin
            _T_185 <= _T_17;
          end else begin
            _T_185 <= 6'h0;
          end
        end else begin
          _T_185 <= _T_187;
        end
      end
    end
    if (reset) begin
      _T_21 <= 6'h0;
    end else begin
      if (_T_12) begin
        if (_T_24) begin
          if (_T_19) begin
            _T_21 <= _T_17;
          end else begin
            _T_21 <= 6'h0;
          end
        end else begin
          _T_21 <= _T_23;
        end
      end
    end
    if (reset) begin
      _T_60 <= 6'h0;
    end else begin
      if (_T_52) begin
        if (_T_63) begin
          if (_T_58) begin
            _T_60 <= _T_57;
          end else begin
            _T_60 <= 6'h0;
          end
        end else begin
          _T_60 <= _T_62;
        end
      end
    end
    if (reset) begin
      _T_79 <= 6'h0;
    end else begin
      if (_T_71) begin
        if (_T_82) begin
          if (_T_77) begin
            _T_79 <= _T_76;
          end else begin
            _T_79 <= 6'h0;
          end
        end else begin
          _T_79 <= _T_81;
        end
      end
    end
  end
endmodule
module dual_ParitalExtractor_1( 
  input        clock, 
  input        reset, 
  input        io_last, 
  output       io_i_ready, 
  input        io_i_valid, 
  input  [2:0] io_i_bits_opcode, 
  output       io_o_valid 
);
  reg [3:0] state; 
  reg [31:0] _RAND_0;
  wire  enable; 
  wire  empty; 
  wire  _GEN_1; 
  wire  _T_19; 
  wire [3:0] _T_23; 
  assign enable = io_i_bits_opcode == 3'h1; 
  assign empty = state == 4'h0; 
  assign _GEN_1 = empty ? 1'h0 : io_i_valid; 
  assign _T_19 = io_i_ready & io_i_valid; 
  assign _T_23 = state - 4'h1; 
  assign io_i_ready = 1'h1; 
  assign io_o_valid = enable ? _GEN_1 : io_i_valid; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      state <= 4'h0;
    end else begin
      if (enable) begin
        if (_T_19) begin
          if (io_last) begin
            state <= 4'h0;
          end else begin
            if (empty) begin
              state <= 4'h8;
            end else begin
              state <= _T_23;
            end
          end
        end
      end
    end
  end
endmodule
module dual_ParitalExtractor( 
  input         clock, 
  input         reset, 
  input         io_last, 
  output        io_i_ready, 
  input         io_i_valid, 
  input  [2:0]  io_i_bits_opcode, 
  input  [2:0]  io_i_bits_param, 
  input  [3:0]  io_i_bits_size, 
  input  [5:0]  io_i_bits_source, 
  input  [31:0] io_i_bits_address, 
  input  [3:0]  io_i_bits_mask, 
  input  [31:0] io_i_bits_data, 
  input         io_o_ready, 
  output        io_o_valid, 
  output [2:0]  io_o_bits_opcode, 
  output [2:0]  io_o_bits_param, 
  output [3:0]  io_o_bits_size, 
  output [5:0]  io_o_bits_source, 
  output [31:0] io_o_bits_address, 
  output [3:0]  io_o_bits_mask, 
  output [31:0] io_o_bits_data 
);
  reg [3:0] state; 
  reg [31:0] _RAND_0;
  reg [31:0] shift; 
  reg [31:0] _RAND_1;
  wire  enable; 
  wire  empty; 
  wire [5:0] _T; 
  wire [94:0] _GEN_12; 
  wire [94:0] _T_1; 
  wire [94:0] _GEN_13; 
  wire [94:0] _T_2; 
  wire [7:0] _T_3; 
  wire [7:0] _T_4; 
  wire [7:0] _T_5; 
  wire [7:0] _T_6; 
  wire [31:0] _T_10; 
  wire  _T_11; 
  wire  _T_12; 
  wire  _T_13; 
  wire  _T_14; 
  wire [3:0] _T_18; 
  wire  _GEN_0; 
  wire  _GEN_1; 
  wire  _T_19; 
  wire [58:0] _T_20; 
  wire [58:0] _T_21; 
  wire [3:0] _T_23; 
  wire [58:0] _GEN_4; 
  wire [58:0] _GEN_10; 
  assign enable = io_i_bits_opcode == 3'h1; 
  assign empty = state == 4'h0; 
  assign _T = {state, 2'h0}; 
  assign _GEN_12 = {{63'd0}, io_i_bits_data}; 
  assign _T_1 = _GEN_12 << _T; 
  assign _GEN_13 = {{63'd0}, shift}; 
  assign _T_2 = _GEN_13 | _T_1; 
  assign _T_3 = _T_2[8:1]; 
  assign _T_4 = _T_2[17:10]; 
  assign _T_5 = _T_2[26:19]; 
  assign _T_6 = _T_2[35:28]; 
  assign _T_10 = {_T_6,_T_5,_T_4,_T_3}; 
  assign _T_11 = _T_2[0]; 
  assign _T_12 = _T_2[9]; 
  assign _T_13 = _T_2[18]; 
  assign _T_14 = _T_2[27]; 
  assign _T_18 = {_T_14,_T_13,_T_12,_T_11}; 
  assign _GEN_0 = empty ? 1'h1 : io_o_ready; 
  assign _GEN_1 = empty ? 1'h0 : io_i_valid; 
  assign _T_19 = io_i_ready & io_i_valid; 
  assign _T_20 = _T_2[94:36]; 
  assign _T_21 = empty ? {{27'd0}, io_i_bits_data} : _T_20; 
  assign _T_23 = state - 4'h1; 
  assign _GEN_4 = _T_19 ? _T_21 : {{27'd0}, shift}; 
  assign _GEN_10 = enable ? _GEN_4 : {{27'd0}, shift}; 
  assign io_i_ready = enable ? _GEN_0 : io_o_ready; 
  assign io_o_valid = enable ? _GEN_1 : io_i_valid; 
  assign io_o_bits_opcode = io_i_bits_opcode; 
  assign io_o_bits_param = io_i_bits_param; 
  assign io_o_bits_size = io_i_bits_size; 
  assign io_o_bits_source = io_i_bits_source; 
  assign io_o_bits_address = io_i_bits_address; 
  assign io_o_bits_mask = enable ? _T_18 : io_i_bits_mask; 
  assign io_o_bits_data = enable ? _T_10 : io_i_bits_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  shift = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      state <= 4'h0;
    end else begin
      if (enable) begin
        if (_T_19) begin
          if (io_last) begin
            state <= 4'h0;
          end else begin
            if (empty) begin
              state <= 4'h8;
            end else begin
              state <= _T_23;
            end
          end
        end
      end
    end
    shift <= _GEN_10[31:0];
  end
endmodule
module dual_PartialInjector( 
  input         clock, 
  input         reset, 
  input         io_i_last, 
  output        io_o_last, 
  output        io_i_ready, 
  input         io_i_valid, 
  input  [2:0]  io_i_bits_opcode, 
  input  [2:0]  io_i_bits_param, 
  input  [2:0]  io_i_bits_size, 
  input  [2:0]  io_i_bits_source, 
  input  [31:0] io_i_bits_address, 
  input  [3:0]  io_i_bits_mask, 
  input  [31:0] io_i_bits_data, 
  input         io_o_ready, 
  output        io_o_valid, 
  output [2:0]  io_o_bits_opcode, 
  output [2:0]  io_o_bits_param, 
  output [2:0]  io_o_bits_size, 
  output [2:0]  io_o_bits_source, 
  output [31:0] io_o_bits_address, 
  output [31:0] io_o_bits_data 
);
  reg [3:0] state; 
  reg [31:0] _RAND_0;
  reg [31:0] shift; 
  reg [31:0] _RAND_1;
  wire  full; 
  wire  partial; 
  reg  last; 
  reg [31:0] _RAND_2;
  wire [7:0] _T_1; 
  wire [7:0] _T_2; 
  wire [7:0] _T_3; 
  wire [7:0] _T_4; 
  wire  _T_5; 
  wire  _T_6; 
  wire  _T_7; 
  wire  _T_8; 
  wire [35:0] _T_15; 
  wire [5:0] _T_16; 
  wire [98:0] _GEN_11; 
  wire [98:0] _T_17; 
  wire [98:0] _GEN_12; 
  wire [98:0] _T_18; 
  wire  _T_19; 
  wire  _T_20; 
  wire  _T_21; 
  wire  _GEN_0; 
  wire  _T_22; 
  wire [66:0] _T_23; 
  wire [3:0] _T_25; 
  wire  _T_26; 
  wire [66:0] _GEN_2; 
  wire  _T_28; 
  wire [66:0] _GEN_3; 
  wire [98:0] _GEN_6; 
  wire [66:0] _GEN_8; 
  assign full = state[3]; 
  assign partial = io_i_bits_opcode == 3'h1; 
  assign _T_1 = io_i_bits_data[7:0]; 
  assign _T_2 = io_i_bits_data[15:8]; 
  assign _T_3 = io_i_bits_data[23:16]; 
  assign _T_4 = io_i_bits_data[31:24]; 
  assign _T_5 = io_i_bits_mask[0]; 
  assign _T_6 = io_i_bits_mask[1]; 
  assign _T_7 = io_i_bits_mask[2]; 
  assign _T_8 = io_i_bits_mask[3]; 
  assign _T_15 = {_T_4,_T_8,_T_3,_T_7,_T_2,_T_6,_T_1,_T_5}; 
  assign _T_16 = {state, 2'h0}; 
  assign _GEN_11 = {{63'd0}, _T_15}; 
  assign _T_17 = _GEN_11 << _T_16; 
  assign _GEN_12 = {{67'd0}, shift}; 
  assign _T_18 = _GEN_12 | _T_17; 
  assign _T_19 = io_i_last | full; 
  assign _T_20 = last == 1'h0; 
  assign _T_21 = _T_19 & _T_20; 
  assign _GEN_0 = _T_21 ? 1'h0 : io_o_ready; 
  assign _T_22 = io_o_ready & io_o_valid; 
  assign _T_23 = _T_18[98:32]; 
  assign _T_25 = state + 4'h1; 
  assign _T_26 = full | last; 
  assign _GEN_2 = _T_26 ? 67'h0 : _T_23; 
  assign _T_28 = io_i_last & _T_20; 
  assign _GEN_3 = _T_22 ? _GEN_2 : {{35'd0}, shift}; 
  assign _GEN_6 = partial ? _T_18 : {{67'd0}, io_i_bits_data}; 
  assign _GEN_8 = partial ? _GEN_3 : {{35'd0}, shift}; 
  assign io_o_last = partial ? last : io_i_last; 
  assign io_i_ready = partial ? _GEN_0 : io_o_ready; 
  assign io_o_valid = io_i_valid; 
  assign io_o_bits_opcode = io_i_bits_opcode; 
  assign io_o_bits_param = io_i_bits_param; 
  assign io_o_bits_size = io_i_bits_size; 
  assign io_o_bits_source = io_i_bits_source; 
  assign io_o_bits_address = io_i_bits_address; 
  assign io_o_bits_data = _GEN_6[31:0]; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  shift = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  last = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      state <= 4'h0;
    end else begin
      if (partial) begin
        if (_T_22) begin
          if (_T_26) begin
            state <= 4'h0;
          end else begin
            state <= _T_25;
          end
        end
      end
    end
    if (reset) begin
      shift <= 32'h0;
    end else begin
      shift <= _GEN_8[31:0];
    end
    if (reset) begin
      last <= 1'h0;
    end else begin
      if (partial) begin
        if (_T_22) begin
          last <= _T_28;
        end
      end
    end
  end
endmodule
module dual_plusarg_reader #(parameter FORMAT="borked=%d", DEFAULT=0) (
   output [31:0] out
);

`ifdef SYNTHESIS
assign out = DEFAULT;
`else
reg [31:0] myplus;
assign out = myplus;

initial begin
   if (!$value$plusargs(FORMAT, myplus)) myplus = DEFAULT;
end
`endif

endmodule
module dual_Queue_14( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [11:0] io_enq_bits, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [11:0] io_deq_bits 
);
  reg [11:0] _T [0:16]; 
  reg [31:0] _RAND_0;
  wire [11:0] _T__T_18_data; 
  wire [4:0] _T__T_18_addr; 
  reg [31:0] _RAND_1;
  wire [11:0] _T__T_10_data; 
  wire [4:0] _T__T_10_addr; 
  wire  _T__T_10_mask; 
  wire  _T__T_10_en; 
  reg [4:0] value; 
  reg [31:0] _RAND_2;
  reg [4:0] value_1; 
  reg [31:0] _RAND_3;
  reg  _T_1; 
  reg [31:0] _RAND_4;
  wire  _T_2; 
  wire  _T_3; 
  wire  _T_4; 
  wire  _T_5; 
  wire  _T_6; 
  wire  _T_8; 
  wire  wrap; 
  wire [4:0] _T_12; 
  wire  wrap_1; 
  wire [4:0] _T_14; 
  wire  _T_15; 
  assign _T__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__T_18_data = _T[_T__T_18_addr]; 
  `else
  assign _T__T_18_data = _T__T_18_addr >= 5'h11 ? _RAND_1[11:0] : _T[_T__T_18_addr]; 
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = value;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; 
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_4 = _T_2 & _T_3; 
  assign _T_5 = _T_2 & _T_1; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign wrap = value == 5'h10; 
  assign _T_12 = value + 5'h1; 
  assign wrap_1 = value_1 == 5'h10; 
  assign _T_14 = value_1 + 5'h1; 
  assign _T_15 = _T_6 != _T_8; 
  assign io_enq_ready = _T_5 == 1'h0; 
  assign io_deq_valid = _T_4 == 1'h0; 
  assign io_deq_bits = _T__T_18_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 17; initvar = initvar+1)
    _T[initvar] = _RAND_0[11:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; 
    end
    if (reset) begin
      value <= 5'h0;
    end else begin
      if (_T_6) begin
        if (wrap) begin
          value <= 5'h0;
        end else begin
          value <= _T_12;
        end
      end
    end
    if (reset) begin
      value_1 <= 5'h0;
    end else begin
      if (_T_8) begin
        if (wrap_1) begin
          value_1 <= 5'h0;
        end else begin
          value_1 <= _T_14;
        end
      end
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_15) begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module dual_Queue_21( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [11:0] io_enq_bits, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [11:0] io_deq_bits 
);
  reg [11:0] _T [0:0]; 
  reg [31:0] _RAND_0;
  wire [11:0] _T__T_14_data; 
  wire  _T__T_14_addr; 
  wire [11:0] _T__T_10_data; 
  wire  _T__T_10_addr; 
  wire  _T__T_10_mask; 
  wire  _T__T_10_en; 
  reg  _T_1; 
  reg [31:0] _RAND_1;
  wire  _T_3; 
  wire  _T_6; 
  wire  _T_8; 
  wire  _T_11; 
  assign _T__T_14_addr = 1'h0;
  assign _T__T_14_data = _T[_T__T_14_addr]; 
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = 1'h0;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _T_11 = _T_6 != _T_8; 
  assign io_enq_ready = _T_1 == 1'h0; 
  assign io_deq_valid = _T_3 == 1'h0; 
  assign io_deq_bits = _T__T_14_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T[initvar] = _RAND_0[11:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; 
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_11) begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module dual_Queue_2( 
  input        clock, 
  input        reset, 
  output       io_enq_ready, 
  input        io_enq_valid, 
  input  [2:0] io_enq_bits_opcode, 
  input  [3:0] io_enq_bits_size, 
  input  [2:0] io_enq_bits_source, 
  input        io_deq_ready, 
  output       io_deq_valid, 
  output [2:0] io_deq_bits_opcode, 
  output [3:0] io_deq_bits_size, 
  output [2:0] io_deq_bits_source 
);
  reg [2:0] _T_opcode [0:0]; 
  reg [31:0] _RAND_0;
  wire [2:0] _T_opcode__T_14_data; 
  wire  _T_opcode__T_14_addr; 
  wire [2:0] _T_opcode__T_10_data; 
  wire  _T_opcode__T_10_addr; 
  wire  _T_opcode__T_10_mask; 
  wire  _T_opcode__T_10_en; 
  reg [3:0] _T_size [0:0]; 
  reg [31:0] _RAND_1;
  wire [3:0] _T_size__T_14_data; 
  wire  _T_size__T_14_addr; 
  wire [3:0] _T_size__T_10_data; 
  wire  _T_size__T_10_addr; 
  wire  _T_size__T_10_mask; 
  wire  _T_size__T_10_en; 
  reg [2:0] _T_source [0:0]; 
  reg [31:0] _RAND_2;
  wire [2:0] _T_source__T_14_data; 
  wire  _T_source__T_14_addr; 
  wire [2:0] _T_source__T_10_data; 
  wire  _T_source__T_10_addr; 
  wire  _T_source__T_10_mask; 
  wire  _T_source__T_10_en; 
  reg  _T_1; 
  reg [31:0] _RAND_3;
  wire  _T_3; 
  wire  _T_6; 
  wire  _T_8; 
  wire  _T_11; 
  assign _T_opcode__T_14_addr = 1'h0;
  assign _T_opcode__T_14_data = _T_opcode[_T_opcode__T_14_addr]; 
  assign _T_opcode__T_10_data = io_enq_bits_opcode;
  assign _T_opcode__T_10_addr = 1'h0;
  assign _T_opcode__T_10_mask = 1'h1;
  assign _T_opcode__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_size__T_14_addr = 1'h0;
  assign _T_size__T_14_data = _T_size[_T_size__T_14_addr]; 
  assign _T_size__T_10_data = io_enq_bits_size;
  assign _T_size__T_10_addr = 1'h0;
  assign _T_size__T_10_mask = 1'h1;
  assign _T_size__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_source__T_14_addr = 1'h0;
  assign _T_source__T_14_data = _T_source[_T_source__T_14_addr]; 
  assign _T_source__T_10_data = io_enq_bits_source;
  assign _T_source__T_10_addr = 1'h0;
  assign _T_source__T_10_mask = 1'h1;
  assign _T_source__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _T_11 = _T_6 != _T_8; 
  assign io_enq_ready = _T_1 == 1'h0; 
  assign io_deq_valid = _T_3 == 1'h0; 
  assign io_deq_bits_opcode = _T_opcode__T_14_data; 
  assign io_deq_bits_size = _T_size__T_14_data; 
  assign io_deq_bits_source = _T_source__T_14_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_size[initvar] = _RAND_1[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_source[initvar] = _RAND_2[2:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T_opcode__T_10_en & _T_opcode__T_10_mask) begin
      _T_opcode[_T_opcode__T_10_addr] <= _T_opcode__T_10_data; 
    end
    if(_T_size__T_10_en & _T_size__T_10_mask) begin
      _T_size[_T_size__T_10_addr] <= _T_size__T_10_data; 
    end
    if(_T_source__T_10_en & _T_source__T_10_mask) begin
      _T_source[_T_source__T_10_addr] <= _T_source__T_10_data; 
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_11) begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module dual_Queue_46( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [63:0] io_enq_bits_data, 
  input  [7:0]  io_enq_bits_strb, 
  input         io_enq_bits_last, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [63:0] io_deq_bits_data, 
  output [7:0]  io_deq_bits_strb, 
  output        io_deq_bits_last 
);
  reg [63:0] _T_data [0:0]; 
  reg [63:0] _RAND_0;
  wire [63:0] _T_data__T_14_data; 
  wire  _T_data__T_14_addr; 
  wire [63:0] _T_data__T_10_data; 
  wire  _T_data__T_10_addr; 
  wire  _T_data__T_10_mask; 
  wire  _T_data__T_10_en; 
  reg [7:0] _T_strb [0:0]; 
  reg [31:0] _RAND_1;
  wire [7:0] _T_strb__T_14_data; 
  wire  _T_strb__T_14_addr; 
  wire [7:0] _T_strb__T_10_data; 
  wire  _T_strb__T_10_addr; 
  wire  _T_strb__T_10_mask; 
  wire  _T_strb__T_10_en; 
  reg  _T_last [0:0]; 
  reg [31:0] _RAND_2;
  wire  _T_last__T_14_data; 
  wire  _T_last__T_14_addr; 
  wire  _T_last__T_10_data; 
  wire  _T_last__T_10_addr; 
  wire  _T_last__T_10_mask; 
  wire  _T_last__T_10_en; 
  reg  _T_1; 
  reg [31:0] _RAND_3;
  wire  _T_3; 
  wire  _T_6; 
  wire  _T_8; 
  wire  _GEN_9; 
  wire  _GEN_14; 
  wire  _GEN_13; 
  wire  _T_11; 
  wire  _T_12; 
  assign _T_data__T_14_addr = 1'h0;
  assign _T_data__T_14_data = _T_data[_T_data__T_14_addr]; 
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = 1'h0;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = _T_3 ? _GEN_9 : _T_6;
  assign _T_strb__T_14_addr = 1'h0;
  assign _T_strb__T_14_data = _T_strb[_T_strb__T_14_addr]; 
  assign _T_strb__T_10_data = io_enq_bits_strb;
  assign _T_strb__T_10_addr = 1'h0;
  assign _T_strb__T_10_mask = 1'h1;
  assign _T_strb__T_10_en = _T_3 ? _GEN_9 : _T_6;
  assign _T_last__T_14_addr = 1'h0;
  assign _T_last__T_14_data = _T_last[_T_last__T_14_addr]; 
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = 1'h0;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = _T_3 ? _GEN_9 : _T_6;
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _GEN_9 = io_deq_ready ? 1'h0 : _T_6; 
  assign _GEN_14 = _T_3 ? _GEN_9 : _T_6; 
  assign _GEN_13 = _T_3 ? 1'h0 : _T_8; 
  assign _T_11 = _GEN_14 != _GEN_13; 
  assign _T_12 = _T_3 == 1'h0; 
  assign io_enq_ready = _T_1 == 1'h0; 
  assign io_deq_valid = io_enq_valid ? 1'h1 : _T_12; 
  assign io_deq_bits_data = _T_3 ? io_enq_bits_data : _T_data__T_14_data; 
  assign io_deq_bits_strb = _T_3 ? io_enq_bits_strb : _T_strb__T_14_data; 
  assign io_deq_bits_last = _T_3 ? io_enq_bits_last : _T_last__T_14_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_strb[initvar] = _RAND_1[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_last[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; 
    end
    if(_T_strb__T_10_en & _T_strb__T_10_mask) begin
      _T_strb[_T_strb__T_10_addr] <= _T_strb__T_10_data; 
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; 
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_3) begin
          if (io_deq_ready) begin
            _T_1 <= 1'h0;
          end else begin
            _T_1 <= _T_6;
          end
        end else begin
          _T_1 <= _T_6;
        end
      end
    end
  end
endmodule
module dual_Queue_47( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [4:0]  io_enq_bits_id, 
  input  [31:0] io_enq_bits_addr, 
  input  [7:0]  io_enq_bits_len, 
  input  [2:0]  io_enq_bits_size, 
  input  [10:0] io_enq_bits_user, 
  input         io_enq_bits_wen, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [4:0]  io_deq_bits_id, 
  output [31:0] io_deq_bits_addr, 
  output [7:0]  io_deq_bits_len, 
  output [2:0]  io_deq_bits_size, 
  output [1:0]  io_deq_bits_burst, 
  output        io_deq_bits_lock, 
  output [3:0]  io_deq_bits_cache, 
  output [2:0]  io_deq_bits_prot, 
  output [3:0]  io_deq_bits_qos, 
  output [10:0] io_deq_bits_user, 
  output [63:0] io_deq_bits_instret, 
  output        io_deq_bits_wen 
);
  reg [4:0] _T_id [0:0]; 
  reg [31:0] _RAND_0;
  wire [4:0] _T_id__T_14_data; 
  wire  _T_id__T_14_addr; 
  wire [4:0] _T_id__T_10_data; 
  wire  _T_id__T_10_addr; 
  wire  _T_id__T_10_mask; 
  wire  _T_id__T_10_en; 
  reg [31:0] _T_addr [0:0]; 
  reg [31:0] _RAND_1;
  wire [31:0] _T_addr__T_14_data; 
  wire  _T_addr__T_14_addr; 
  wire [31:0] _T_addr__T_10_data; 
  wire  _T_addr__T_10_addr; 
  wire  _T_addr__T_10_mask; 
  wire  _T_addr__T_10_en; 
  reg [7:0] _T_len [0:0]; 
  reg [31:0] _RAND_2;
  wire [7:0] _T_len__T_14_data; 
  wire  _T_len__T_14_addr; 
  wire [7:0] _T_len__T_10_data; 
  wire  _T_len__T_10_addr; 
  wire  _T_len__T_10_mask; 
  wire  _T_len__T_10_en; 
  reg [2:0] _T_size [0:0]; 
  reg [31:0] _RAND_3;
  wire [2:0] _T_size__T_14_data; 
  wire  _T_size__T_14_addr; 
  wire [2:0] _T_size__T_10_data; 
  wire  _T_size__T_10_addr; 
  wire  _T_size__T_10_mask; 
  wire  _T_size__T_10_en; 
  reg [1:0] _T_burst [0:0]; 
  reg [31:0] _RAND_4;
  wire [1:0] _T_burst__T_14_data; 
  wire  _T_burst__T_14_addr; 
  wire [1:0] _T_burst__T_10_data; 
  wire  _T_burst__T_10_addr; 
  wire  _T_burst__T_10_mask; 
  wire  _T_burst__T_10_en; 
  reg  _T_lock [0:0]; 
  reg [31:0] _RAND_5;
  wire  _T_lock__T_14_data; 
  wire  _T_lock__T_14_addr; 
  wire  _T_lock__T_10_data; 
  wire  _T_lock__T_10_addr; 
  wire  _T_lock__T_10_mask; 
  wire  _T_lock__T_10_en; 
  reg [3:0] _T_cache [0:0]; 
  reg [31:0] _RAND_6;
  wire [3:0] _T_cache__T_14_data; 
  wire  _T_cache__T_14_addr; 
  wire [3:0] _T_cache__T_10_data; 
  wire  _T_cache__T_10_addr; 
  wire  _T_cache__T_10_mask; 
  wire  _T_cache__T_10_en; 
  reg [2:0] _T_prot [0:0]; 
  reg [31:0] _RAND_7;
  wire [2:0] _T_prot__T_14_data; 
  wire  _T_prot__T_14_addr; 
  wire [2:0] _T_prot__T_10_data; 
  wire  _T_prot__T_10_addr; 
  wire  _T_prot__T_10_mask; 
  wire  _T_prot__T_10_en; 
  reg [3:0] _T_qos [0:0]; 
  reg [31:0] _RAND_8;
  wire [3:0] _T_qos__T_14_data; 
  wire  _T_qos__T_14_addr; 
  wire [3:0] _T_qos__T_10_data; 
  wire  _T_qos__T_10_addr; 
  wire  _T_qos__T_10_mask; 
  wire  _T_qos__T_10_en; 
  reg [10:0] _T_user [0:0]; 
  reg [31:0] _RAND_9;
  wire [10:0] _T_user__T_14_data; 
  wire  _T_user__T_14_addr; 
  wire [10:0] _T_user__T_10_data; 
  wire  _T_user__T_10_addr; 
  wire  _T_user__T_10_mask; 
  wire  _T_user__T_10_en; 
  reg [63:0] _T_instret [0:0]; 
  reg [63:0] _RAND_10;
  wire [63:0] _T_instret__T_14_data; 
  wire  _T_instret__T_14_addr; 
  wire [63:0] _T_instret__T_10_data; 
  wire  _T_instret__T_10_addr; 
  wire  _T_instret__T_10_mask; 
  wire  _T_instret__T_10_en; 
  reg  _T_wen [0:0]; 
  reg [31:0] _RAND_11;
  wire  _T_wen__T_14_data; 
  wire  _T_wen__T_14_addr; 
  wire  _T_wen__T_10_data; 
  wire  _T_wen__T_10_addr; 
  wire  _T_wen__T_10_mask; 
  wire  _T_wen__T_10_en; 
  reg  _T_1; 
  reg [31:0] _RAND_12;
  wire  _T_3; 
  wire  _T_6; 
  wire  _T_8; 
  wire  _GEN_18; 
  wire  _GEN_32; 
  wire  _GEN_31; 
  wire  _T_11; 
  wire  _T_12; 
  assign _T_id__T_14_addr = 1'h0;
  assign _T_id__T_14_data = _T_id[_T_id__T_14_addr]; 
  assign _T_id__T_10_data = io_enq_bits_id;
  assign _T_id__T_10_addr = 1'h0;
  assign _T_id__T_10_mask = 1'h1;
  assign _T_id__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_addr__T_14_addr = 1'h0;
  assign _T_addr__T_14_data = _T_addr[_T_addr__T_14_addr]; 
  assign _T_addr__T_10_data = io_enq_bits_addr;
  assign _T_addr__T_10_addr = 1'h0;
  assign _T_addr__T_10_mask = 1'h1;
  assign _T_addr__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_len__T_14_addr = 1'h0;
  assign _T_len__T_14_data = _T_len[_T_len__T_14_addr]; 
  assign _T_len__T_10_data = io_enq_bits_len;
  assign _T_len__T_10_addr = 1'h0;
  assign _T_len__T_10_mask = 1'h1;
  assign _T_len__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_size__T_14_addr = 1'h0;
  assign _T_size__T_14_data = _T_size[_T_size__T_14_addr]; 
  assign _T_size__T_10_data = io_enq_bits_size;
  assign _T_size__T_10_addr = 1'h0;
  assign _T_size__T_10_mask = 1'h1;
  assign _T_size__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_burst__T_14_addr = 1'h0;
  assign _T_burst__T_14_data = _T_burst[_T_burst__T_14_addr]; 
  assign _T_burst__T_10_data = 2'h1;
  assign _T_burst__T_10_addr = 1'h0;
  assign _T_burst__T_10_mask = 1'h1;
  assign _T_burst__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_lock__T_14_addr = 1'h0;
  assign _T_lock__T_14_data = _T_lock[_T_lock__T_14_addr]; 
  assign _T_lock__T_10_data = 1'h0;
  assign _T_lock__T_10_addr = 1'h0;
  assign _T_lock__T_10_mask = 1'h1;
  assign _T_lock__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_cache__T_14_addr = 1'h0;
  assign _T_cache__T_14_data = _T_cache[_T_cache__T_14_addr]; 
  assign _T_cache__T_10_data = 4'h0;
  assign _T_cache__T_10_addr = 1'h0;
  assign _T_cache__T_10_mask = 1'h1;
  assign _T_cache__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_prot__T_14_addr = 1'h0;
  assign _T_prot__T_14_data = _T_prot[_T_prot__T_14_addr]; 
  assign _T_prot__T_10_data = 3'h1;
  assign _T_prot__T_10_addr = 1'h0;
  assign _T_prot__T_10_mask = 1'h1;
  assign _T_prot__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_qos__T_14_addr = 1'h0;
  assign _T_qos__T_14_data = _T_qos[_T_qos__T_14_addr]; 
  assign _T_qos__T_10_data = 4'h0;
  assign _T_qos__T_10_addr = 1'h0;
  assign _T_qos__T_10_mask = 1'h1;
  assign _T_qos__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_user__T_14_addr = 1'h0;
  assign _T_user__T_14_data = _T_user[_T_user__T_14_addr]; 
  assign _T_user__T_10_data = io_enq_bits_user;
  assign _T_user__T_10_addr = 1'h0;
  assign _T_user__T_10_mask = 1'h1;
  assign _T_user__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_instret__T_14_addr = 1'h0;
  assign _T_instret__T_14_data = _T_instret[_T_instret__T_14_addr]; 
  assign _T_instret__T_10_data = 64'h0;
  assign _T_instret__T_10_addr = 1'h0;
  assign _T_instret__T_10_mask = 1'h1;
  assign _T_instret__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_wen__T_14_addr = 1'h0;
  assign _T_wen__T_14_data = _T_wen[_T_wen__T_14_addr]; 
  assign _T_wen__T_10_data = io_enq_bits_wen;
  assign _T_wen__T_10_addr = 1'h0;
  assign _T_wen__T_10_mask = 1'h1;
  assign _T_wen__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _GEN_18 = io_deq_ready ? 1'h0 : _T_6; 
  assign _GEN_32 = _T_3 ? _GEN_18 : _T_6; 
  assign _GEN_31 = _T_3 ? 1'h0 : _T_8; 
  assign _T_11 = _GEN_32 != _GEN_31; 
  assign _T_12 = _T_3 == 1'h0; 
  assign io_enq_ready = _T_1 == 1'h0; 
  assign io_deq_valid = io_enq_valid ? 1'h1 : _T_12; 
  assign io_deq_bits_id = _T_3 ? io_enq_bits_id : _T_id__T_14_data; 
  assign io_deq_bits_addr = _T_3 ? io_enq_bits_addr : _T_addr__T_14_data; 
  assign io_deq_bits_len = _T_3 ? io_enq_bits_len : _T_len__T_14_data; 
  assign io_deq_bits_size = _T_3 ? io_enq_bits_size : _T_size__T_14_data; 
  assign io_deq_bits_burst = _T_3 ? 2'h1 : _T_burst__T_14_data; 
  assign io_deq_bits_lock = _T_3 ? 1'h0 : _T_lock__T_14_data; 
  assign io_deq_bits_cache = _T_3 ? 4'h0 : _T_cache__T_14_data; 
  assign io_deq_bits_prot = _T_3 ? 3'h1 : _T_prot__T_14_data; 
  assign io_deq_bits_qos = _T_3 ? 4'h0 : _T_qos__T_14_data; 
  assign io_deq_bits_user = _T_3 ? io_enq_bits_user : _T_user__T_14_data; 
  assign io_deq_bits_instret = _T_3 ? 64'h0 : _T_instret__T_14_data; 
  assign io_deq_bits_wen = _T_3 ? io_enq_bits_wen : _T_wen__T_14_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_id[initvar] = _RAND_0[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_addr[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_len[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_size[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_burst[initvar] = _RAND_4[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_lock[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_cache[initvar] = _RAND_6[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_prot[initvar] = _RAND_7[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_qos[initvar] = _RAND_8[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_user[initvar] = _RAND_9[10:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_10 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_instret[initvar] = _RAND_10[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_11 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_wen[initvar] = _RAND_11[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_1 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T_id__T_10_en & _T_id__T_10_mask) begin
      _T_id[_T_id__T_10_addr] <= _T_id__T_10_data; 
    end
    if(_T_addr__T_10_en & _T_addr__T_10_mask) begin
      _T_addr[_T_addr__T_10_addr] <= _T_addr__T_10_data; 
    end
    if(_T_len__T_10_en & _T_len__T_10_mask) begin
      _T_len[_T_len__T_10_addr] <= _T_len__T_10_data; 
    end
    if(_T_size__T_10_en & _T_size__T_10_mask) begin
      _T_size[_T_size__T_10_addr] <= _T_size__T_10_data; 
    end
    if(_T_burst__T_10_en & _T_burst__T_10_mask) begin
      _T_burst[_T_burst__T_10_addr] <= _T_burst__T_10_data; 
    end
    if(_T_lock__T_10_en & _T_lock__T_10_mask) begin
      _T_lock[_T_lock__T_10_addr] <= _T_lock__T_10_data; 
    end
    if(_T_cache__T_10_en & _T_cache__T_10_mask) begin
      _T_cache[_T_cache__T_10_addr] <= _T_cache__T_10_data; 
    end
    if(_T_prot__T_10_en & _T_prot__T_10_mask) begin
      _T_prot[_T_prot__T_10_addr] <= _T_prot__T_10_data; 
    end
    if(_T_qos__T_10_en & _T_qos__T_10_mask) begin
      _T_qos[_T_qos__T_10_addr] <= _T_qos__T_10_data; 
    end
    if(_T_user__T_10_en & _T_user__T_10_mask) begin
      _T_user[_T_user__T_10_addr] <= _T_user__T_10_data; 
    end
    if(_T_instret__T_10_en & _T_instret__T_10_mask) begin
      _T_instret[_T_instret__T_10_addr] <= _T_instret__T_10_data; 
    end
    if(_T_wen__T_10_en & _T_wen__T_10_mask) begin
      _T_wen[_T_wen__T_10_addr] <= _T_wen__T_10_data; 
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_3) begin
          if (io_deq_ready) begin
            _T_1 <= 1'h0;
          end else begin
            _T_1 <= _T_6;
          end
        end else begin
          _T_1 <= _T_6;
        end
      end
    end
  end
endmodule
module dual_Queue_48( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [30:0] io_enq_bits_addr, 
  input  [7:0]  io_enq_bits_len, 
  input  [2:0]  io_enq_bits_size, 
  input  [1:0]  io_enq_bits_burst, 
  input         io_enq_bits_lock, 
  input  [3:0]  io_enq_bits_cache, 
  input  [2:0]  io_enq_bits_prot, 
  input  [3:0]  io_enq_bits_qos, 
  input  [63:0] io_enq_bits_instret, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output        io_deq_bits_id, 
  output [30:0] io_deq_bits_addr, 
  output [7:0]  io_deq_bits_len, 
  output [2:0]  io_deq_bits_size, 
  output [1:0]  io_deq_bits_burst, 
  output        io_deq_bits_lock, 
  output [3:0]  io_deq_bits_cache, 
  output [2:0]  io_deq_bits_prot, 
  output [3:0]  io_deq_bits_qos, 
  output [63:0] io_deq_bits_instret 
);
  reg  _T_id [0:1]; 
  reg [31:0] _RAND_0;
  wire  _T_id__T_18_data; 
  wire  _T_id__T_18_addr; 
  wire  _T_id__T_10_data; 
  wire  _T_id__T_10_addr; 
  wire  _T_id__T_10_mask; 
  wire  _T_id__T_10_en; 
  reg [30:0] _T_addr [0:1]; 
  reg [31:0] _RAND_1;
  wire [30:0] _T_addr__T_18_data; 
  wire  _T_addr__T_18_addr; 
  wire [30:0] _T_addr__T_10_data; 
  wire  _T_addr__T_10_addr; 
  wire  _T_addr__T_10_mask; 
  wire  _T_addr__T_10_en; 
  reg [7:0] _T_len [0:1]; 
  reg [31:0] _RAND_2;
  wire [7:0] _T_len__T_18_data; 
  wire  _T_len__T_18_addr; 
  wire [7:0] _T_len__T_10_data; 
  wire  _T_len__T_10_addr; 
  wire  _T_len__T_10_mask; 
  wire  _T_len__T_10_en; 
  reg [2:0] _T_size [0:1]; 
  reg [31:0] _RAND_3;
  wire [2:0] _T_size__T_18_data; 
  wire  _T_size__T_18_addr; 
  wire [2:0] _T_size__T_10_data; 
  wire  _T_size__T_10_addr; 
  wire  _T_size__T_10_mask; 
  wire  _T_size__T_10_en; 
  reg [1:0] _T_burst [0:1]; 
  reg [31:0] _RAND_4;
  wire [1:0] _T_burst__T_18_data; 
  wire  _T_burst__T_18_addr; 
  wire [1:0] _T_burst__T_10_data; 
  wire  _T_burst__T_10_addr; 
  wire  _T_burst__T_10_mask; 
  wire  _T_burst__T_10_en; 
  reg  _T_lock [0:1]; 
  reg [31:0] _RAND_5;
  wire  _T_lock__T_18_data; 
  wire  _T_lock__T_18_addr; 
  wire  _T_lock__T_10_data; 
  wire  _T_lock__T_10_addr; 
  wire  _T_lock__T_10_mask; 
  wire  _T_lock__T_10_en; 
  reg [3:0] _T_cache [0:1]; 
  reg [31:0] _RAND_6;
  wire [3:0] _T_cache__T_18_data; 
  wire  _T_cache__T_18_addr; 
  wire [3:0] _T_cache__T_10_data; 
  wire  _T_cache__T_10_addr; 
  wire  _T_cache__T_10_mask; 
  wire  _T_cache__T_10_en; 
  reg [2:0] _T_prot [0:1]; 
  reg [31:0] _RAND_7;
  wire [2:0] _T_prot__T_18_data; 
  wire  _T_prot__T_18_addr; 
  wire [2:0] _T_prot__T_10_data; 
  wire  _T_prot__T_10_addr; 
  wire  _T_prot__T_10_mask; 
  wire  _T_prot__T_10_en; 
  reg [3:0] _T_qos [0:1]; 
  reg [31:0] _RAND_8;
  wire [3:0] _T_qos__T_18_data; 
  wire  _T_qos__T_18_addr; 
  wire [3:0] _T_qos__T_10_data; 
  wire  _T_qos__T_10_addr; 
  wire  _T_qos__T_10_mask; 
  wire  _T_qos__T_10_en; 
  reg [63:0] _T_instret [0:1]; 
  reg [63:0] _RAND_9;
  wire [63:0] _T_instret__T_18_data; 
  wire  _T_instret__T_18_addr; 
  wire [63:0] _T_instret__T_10_data; 
  wire  _T_instret__T_10_addr; 
  wire  _T_instret__T_10_mask; 
  wire  _T_instret__T_10_en; 
  reg  value; 
  reg [31:0] _RAND_10;
  reg  value_1; 
  reg [31:0] _RAND_11;
  reg  _T_1; 
  reg [31:0] _RAND_12;
  wire  _T_2; 
  wire  _T_3; 
  wire  _T_4; 
  wire  _T_5; 
  wire  _T_6; 
  wire  _T_8; 
  wire  _T_12; 
  wire  _T_14; 
  wire  _T_15; 
  assign _T_id__T_18_addr = value_1;
  assign _T_id__T_18_data = _T_id[_T_id__T_18_addr]; 
  assign _T_id__T_10_data = 1'h0;
  assign _T_id__T_10_addr = value;
  assign _T_id__T_10_mask = 1'h1;
  assign _T_id__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_addr__T_18_addr = value_1;
  assign _T_addr__T_18_data = _T_addr[_T_addr__T_18_addr]; 
  assign _T_addr__T_10_data = io_enq_bits_addr;
  assign _T_addr__T_10_addr = value;
  assign _T_addr__T_10_mask = 1'h1;
  assign _T_addr__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_len__T_18_addr = value_1;
  assign _T_len__T_18_data = _T_len[_T_len__T_18_addr]; 
  assign _T_len__T_10_data = io_enq_bits_len;
  assign _T_len__T_10_addr = value;
  assign _T_len__T_10_mask = 1'h1;
  assign _T_len__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_size__T_18_addr = value_1;
  assign _T_size__T_18_data = _T_size[_T_size__T_18_addr]; 
  assign _T_size__T_10_data = io_enq_bits_size;
  assign _T_size__T_10_addr = value;
  assign _T_size__T_10_mask = 1'h1;
  assign _T_size__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_burst__T_18_addr = value_1;
  assign _T_burst__T_18_data = _T_burst[_T_burst__T_18_addr]; 
  assign _T_burst__T_10_data = io_enq_bits_burst;
  assign _T_burst__T_10_addr = value;
  assign _T_burst__T_10_mask = 1'h1;
  assign _T_burst__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_lock__T_18_addr = value_1;
  assign _T_lock__T_18_data = _T_lock[_T_lock__T_18_addr]; 
  assign _T_lock__T_10_data = io_enq_bits_lock;
  assign _T_lock__T_10_addr = value;
  assign _T_lock__T_10_mask = 1'h1;
  assign _T_lock__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_cache__T_18_addr = value_1;
  assign _T_cache__T_18_data = _T_cache[_T_cache__T_18_addr]; 
  assign _T_cache__T_10_data = io_enq_bits_cache;
  assign _T_cache__T_10_addr = value;
  assign _T_cache__T_10_mask = 1'h1;
  assign _T_cache__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_prot__T_18_addr = value_1;
  assign _T_prot__T_18_data = _T_prot[_T_prot__T_18_addr]; 
  assign _T_prot__T_10_data = io_enq_bits_prot;
  assign _T_prot__T_10_addr = value;
  assign _T_prot__T_10_mask = 1'h1;
  assign _T_prot__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_qos__T_18_addr = value_1;
  assign _T_qos__T_18_data = _T_qos[_T_qos__T_18_addr]; 
  assign _T_qos__T_10_data = io_enq_bits_qos;
  assign _T_qos__T_10_addr = value;
  assign _T_qos__T_10_mask = 1'h1;
  assign _T_qos__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_instret__T_18_addr = value_1;
  assign _T_instret__T_18_data = _T_instret[_T_instret__T_18_addr]; 
  assign _T_instret__T_10_data = io_enq_bits_instret;
  assign _T_instret__T_10_addr = value;
  assign _T_instret__T_10_mask = 1'h1;
  assign _T_instret__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; 
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_4 = _T_2 & _T_3; 
  assign _T_5 = _T_2 & _T_1; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _T_12 = value + 1'h1; 
  assign _T_14 = value_1 + 1'h1; 
  assign _T_15 = _T_6 != _T_8; 
  assign io_enq_ready = _T_5 == 1'h0; 
  assign io_deq_valid = _T_4 == 1'h0; 
  assign io_deq_bits_id = _T_id__T_18_data; 
  assign io_deq_bits_addr = _T_addr__T_18_data; 
  assign io_deq_bits_len = _T_len__T_18_data; 
  assign io_deq_bits_size = _T_size__T_18_data; 
  assign io_deq_bits_burst = _T_burst__T_18_data; 
  assign io_deq_bits_lock = _T_lock__T_18_data; 
  assign io_deq_bits_cache = _T_cache__T_18_data; 
  assign io_deq_bits_prot = _T_prot__T_18_data; 
  assign io_deq_bits_qos = _T_qos__T_18_data; 
  assign io_deq_bits_instret = _T_instret__T_18_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_id[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_addr[initvar] = _RAND_1[30:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_len[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_size[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_burst[initvar] = _RAND_4[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_lock[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_cache[initvar] = _RAND_6[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_prot[initvar] = _RAND_7[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_qos[initvar] = _RAND_8[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_instret[initvar] = _RAND_9[63:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  value = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  value_1 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_1 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T_id__T_10_en & _T_id__T_10_mask) begin
      _T_id[_T_id__T_10_addr] <= _T_id__T_10_data; 
    end
    if(_T_addr__T_10_en & _T_addr__T_10_mask) begin
      _T_addr[_T_addr__T_10_addr] <= _T_addr__T_10_data; 
    end
    if(_T_len__T_10_en & _T_len__T_10_mask) begin
      _T_len[_T_len__T_10_addr] <= _T_len__T_10_data; 
    end
    if(_T_size__T_10_en & _T_size__T_10_mask) begin
      _T_size[_T_size__T_10_addr] <= _T_size__T_10_data; 
    end
    if(_T_burst__T_10_en & _T_burst__T_10_mask) begin
      _T_burst[_T_burst__T_10_addr] <= _T_burst__T_10_data; 
    end
    if(_T_lock__T_10_en & _T_lock__T_10_mask) begin
      _T_lock[_T_lock__T_10_addr] <= _T_lock__T_10_data; 
    end
    if(_T_cache__T_10_en & _T_cache__T_10_mask) begin
      _T_cache[_T_cache__T_10_addr] <= _T_cache__T_10_data; 
    end
    if(_T_prot__T_10_en & _T_prot__T_10_mask) begin
      _T_prot[_T_prot__T_10_addr] <= _T_prot__T_10_data; 
    end
    if(_T_qos__T_10_en & _T_qos__T_10_mask) begin
      _T_qos[_T_qos__T_10_addr] <= _T_qos__T_10_data; 
    end
    if(_T_instret__T_10_en & _T_instret__T_10_mask) begin
      _T_instret[_T_instret__T_10_addr] <= _T_instret__T_10_data; 
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (_T_6) begin
        value <= _T_12;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (_T_8) begin
        value_1 <= _T_14;
      end
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_15) begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module dual_Queue_49( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [63:0] io_enq_bits_data, 
  input  [7:0]  io_enq_bits_strb, 
  input         io_enq_bits_last, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [63:0] io_deq_bits_data, 
  output [7:0]  io_deq_bits_strb, 
  output        io_deq_bits_last 
);
  reg [63:0] _T_data [0:1]; 
  reg [63:0] _RAND_0;
  wire [63:0] _T_data__T_18_data; 
  wire  _T_data__T_18_addr; 
  wire [63:0] _T_data__T_10_data; 
  wire  _T_data__T_10_addr; 
  wire  _T_data__T_10_mask; 
  wire  _T_data__T_10_en; 
  reg [7:0] _T_strb [0:1]; 
  reg [31:0] _RAND_1;
  wire [7:0] _T_strb__T_18_data; 
  wire  _T_strb__T_18_addr; 
  wire [7:0] _T_strb__T_10_data; 
  wire  _T_strb__T_10_addr; 
  wire  _T_strb__T_10_mask; 
  wire  _T_strb__T_10_en; 
  reg  _T_last [0:1]; 
  reg [31:0] _RAND_2;
  wire  _T_last__T_18_data; 
  wire  _T_last__T_18_addr; 
  wire  _T_last__T_10_data; 
  wire  _T_last__T_10_addr; 
  wire  _T_last__T_10_mask; 
  wire  _T_last__T_10_en; 
  reg  value; 
  reg [31:0] _RAND_3;
  reg  value_1; 
  reg [31:0] _RAND_4;
  reg  _T_1; 
  reg [31:0] _RAND_5;
  wire  _T_2; 
  wire  _T_3; 
  wire  _T_4; 
  wire  _T_5; 
  wire  _T_6; 
  wire  _T_8; 
  wire  _T_12; 
  wire  _T_14; 
  wire  _T_15; 
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; 
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_strb__T_18_addr = value_1;
  assign _T_strb__T_18_data = _T_strb[_T_strb__T_18_addr]; 
  assign _T_strb__T_10_data = io_enq_bits_strb;
  assign _T_strb__T_10_addr = value;
  assign _T_strb__T_10_mask = 1'h1;
  assign _T_strb__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; 
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; 
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_4 = _T_2 & _T_3; 
  assign _T_5 = _T_2 & _T_1; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _T_12 = value + 1'h1; 
  assign _T_14 = value_1 + 1'h1; 
  assign _T_15 = _T_6 != _T_8; 
  assign io_enq_ready = _T_5 == 1'h0; 
  assign io_deq_valid = _T_4 == 1'h0; 
  assign io_deq_bits_data = _T_data__T_18_data; 
  assign io_deq_bits_strb = _T_strb__T_18_data; 
  assign io_deq_bits_last = _T_last__T_18_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_strb[initvar] = _RAND_1[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; 
    end
    if(_T_strb__T_10_en & _T_strb__T_10_mask) begin
      _T_strb[_T_strb__T_10_addr] <= _T_strb__T_10_data; 
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; 
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (_T_6) begin
        value <= _T_12;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (_T_8) begin
        value_1 <= _T_14;
      end
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_15) begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module dual_Queue_4( 
  input         clock, 
  input         reset, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [2:0]  io_deq_bits_opcode, 
  output [2:0]  io_deq_bits_param, 
  output [3:0]  io_deq_bits_size, 
  output        io_deq_bits_source, 
  output [31:0] io_deq_bits_address, 
  output        io_deq_bits_corrupt 
);
  reg [2:0] _T_opcode [0:1]; 
  reg [31:0] _RAND_0;
  wire [2:0] _T_opcode__T_18_data; 
  wire  _T_opcode__T_18_addr; 
  wire [2:0] _T_opcode__T_10_data; 
  wire  _T_opcode__T_10_addr; 
  wire  _T_opcode__T_10_mask; 
  wire  _T_opcode__T_10_en; 
  reg [2:0] _T_param [0:1]; 
  reg [31:0] _RAND_1;
  wire [2:0] _T_param__T_18_data; 
  wire  _T_param__T_18_addr; 
  wire [2:0] _T_param__T_10_data; 
  wire  _T_param__T_10_addr; 
  wire  _T_param__T_10_mask; 
  wire  _T_param__T_10_en; 
  reg [3:0] _T_size [0:1]; 
  reg [31:0] _RAND_2;
  wire [3:0] _T_size__T_18_data; 
  wire  _T_size__T_18_addr; 
  wire [3:0] _T_size__T_10_data; 
  wire  _T_size__T_10_addr; 
  wire  _T_size__T_10_mask; 
  wire  _T_size__T_10_en; 
  reg  _T_source [0:1]; 
  reg [31:0] _RAND_3;
  wire  _T_source__T_18_data; 
  wire  _T_source__T_18_addr; 
  wire  _T_source__T_10_data; 
  wire  _T_source__T_10_addr; 
  wire  _T_source__T_10_mask; 
  wire  _T_source__T_10_en; 
  reg [31:0] _T_address [0:1]; 
  reg [31:0] _RAND_4;
  wire [31:0] _T_address__T_18_data; 
  wire  _T_address__T_18_addr; 
  wire [31:0] _T_address__T_10_data; 
  wire  _T_address__T_10_addr; 
  wire  _T_address__T_10_mask; 
  wire  _T_address__T_10_en; 
  reg  _T_corrupt [0:1]; 
  reg [31:0] _RAND_5;
  wire  _T_corrupt__T_18_data; 
  wire  _T_corrupt__T_18_addr; 
  wire  _T_corrupt__T_10_data; 
  wire  _T_corrupt__T_10_addr; 
  wire  _T_corrupt__T_10_mask; 
  wire  _T_corrupt__T_10_en; 
  reg  value_1; 
  reg [31:0] _RAND_6;
  wire  _T_2; 
  wire  _T_8; 
  wire  _T_14; 
  assign _T_opcode__T_18_addr = value_1;
  assign _T_opcode__T_18_data = _T_opcode[_T_opcode__T_18_addr]; 
  assign _T_opcode__T_10_data = 3'h4;
  assign _T_opcode__T_10_addr = 1'h0;
  assign _T_opcode__T_10_mask = 1'h1;
  assign _T_opcode__T_10_en = 1'h0;
  assign _T_param__T_18_addr = value_1;
  assign _T_param__T_18_data = _T_param[_T_param__T_18_addr]; 
  assign _T_param__T_10_data = 3'h5;
  assign _T_param__T_10_addr = 1'h0;
  assign _T_param__T_10_mask = 1'h1;
  assign _T_param__T_10_en = 1'h0;
  assign _T_size__T_18_addr = value_1;
  assign _T_size__T_18_data = _T_size[_T_size__T_18_addr]; 
  assign _T_size__T_10_data = 4'h0;
  assign _T_size__T_10_addr = 1'h0;
  assign _T_size__T_10_mask = 1'h1;
  assign _T_size__T_10_en = 1'h0;
  assign _T_source__T_18_addr = value_1;
  assign _T_source__T_18_data = _T_source[_T_source__T_18_addr]; 
  assign _T_source__T_10_data = 1'h0;
  assign _T_source__T_10_addr = 1'h0;
  assign _T_source__T_10_mask = 1'h1;
  assign _T_source__T_10_en = 1'h0;
  assign _T_address__T_18_addr = value_1;
  assign _T_address__T_18_data = _T_address[_T_address__T_18_addr]; 
  assign _T_address__T_10_data = 32'h0;
  assign _T_address__T_10_addr = 1'h0;
  assign _T_address__T_10_mask = 1'h1;
  assign _T_address__T_10_en = 1'h0;
  assign _T_corrupt__T_18_addr = value_1;
  assign _T_corrupt__T_18_data = _T_corrupt[_T_corrupt__T_18_addr]; 
  assign _T_corrupt__T_10_data = 1'h0;
  assign _T_corrupt__T_10_addr = 1'h0;
  assign _T_corrupt__T_10_mask = 1'h1;
  assign _T_corrupt__T_10_en = 1'h0;
  assign _T_2 = 1'h0 == value_1; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _T_14 = value_1 + 1'h1; 
  assign io_deq_valid = _T_2 == 1'h0; 
  assign io_deq_bits_opcode = _T_opcode__T_18_data; 
  assign io_deq_bits_param = _T_param__T_18_data; 
  assign io_deq_bits_size = _T_size__T_18_data; 
  assign io_deq_bits_source = _T_source__T_18_data; 
  assign io_deq_bits_address = _T_address__T_18_data; 
  assign io_deq_bits_corrupt = _T_corrupt__T_18_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_param[initvar] = _RAND_1[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_size[initvar] = _RAND_2[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_source[initvar] = _RAND_3[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_address[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_corrupt[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  value_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T_opcode__T_10_en & _T_opcode__T_10_mask) begin
      _T_opcode[_T_opcode__T_10_addr] <= _T_opcode__T_10_data; 
    end
    if(_T_param__T_10_en & _T_param__T_10_mask) begin
      _T_param[_T_param__T_10_addr] <= _T_param__T_10_data; 
    end
    if(_T_size__T_10_en & _T_size__T_10_mask) begin
      _T_size[_T_size__T_10_addr] <= _T_size__T_10_data; 
    end
    if(_T_source__T_10_en & _T_source__T_10_mask) begin
      _T_source[_T_source__T_10_addr] <= _T_source__T_10_data; 
    end
    if(_T_address__T_10_en & _T_address__T_10_mask) begin
      _T_address[_T_address__T_10_addr] <= _T_address__T_10_data; 
    end
    if(_T_corrupt__T_10_en & _T_corrupt__T_10_mask) begin
      _T_corrupt[_T_corrupt__T_10_addr] <= _T_corrupt__T_10_data; 
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (_T_8) begin
        value_1 <= _T_14;
      end
    end
  end
endmodule
module dual_Queue_50( 
  input        clock, 
  input        reset, 
  output       io_enq_ready, 
  input        io_enq_valid, 
  input  [1:0] io_enq_bits_resp, 
  input        io_deq_ready, 
  output       io_deq_valid, 
  output [1:0] io_deq_bits_resp 
);
  reg [1:0] _T_resp [0:1]; 
  reg [31:0] _RAND_0;
  wire [1:0] _T_resp__T_18_data; 
  wire  _T_resp__T_18_addr; 
  wire [1:0] _T_resp__T_10_data; 
  wire  _T_resp__T_10_addr; 
  wire  _T_resp__T_10_mask; 
  wire  _T_resp__T_10_en; 
  reg  value; 
  reg [31:0] _RAND_1;
  reg  value_1; 
  reg [31:0] _RAND_2;
  reg  _T_1; 
  reg [31:0] _RAND_3;
  wire  _T_2; 
  wire  _T_3; 
  wire  _T_4; 
  wire  _T_5; 
  wire  _T_6; 
  wire  _T_8; 
  wire  _T_12; 
  wire  _T_14; 
  wire  _T_15; 
  assign _T_resp__T_18_addr = value_1;
  assign _T_resp__T_18_data = _T_resp[_T_resp__T_18_addr]; 
  assign _T_resp__T_10_data = io_enq_bits_resp;
  assign _T_resp__T_10_addr = value;
  assign _T_resp__T_10_mask = 1'h1;
  assign _T_resp__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; 
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_4 = _T_2 & _T_3; 
  assign _T_5 = _T_2 & _T_1; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _T_12 = value + 1'h1; 
  assign _T_14 = value_1 + 1'h1; 
  assign _T_15 = _T_6 != _T_8; 
  assign io_enq_ready = _T_5 == 1'h0; 
  assign io_deq_valid = _T_4 == 1'h0; 
  assign io_deq_bits_resp = _T_resp__T_18_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_resp[initvar] = _RAND_0[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T_resp__T_10_en & _T_resp__T_10_mask) begin
      _T_resp[_T_resp__T_10_addr] <= _T_resp__T_10_data; 
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (_T_6) begin
        value <= _T_12;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (_T_8) begin
        value_1 <= _T_14;
      end
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_15) begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module dual_Queue_52( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [63:0] io_enq_bits_data, 
  input  [1:0]  io_enq_bits_resp, 
  input         io_enq_bits_last, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [63:0] io_deq_bits_data, 
  output [1:0]  io_deq_bits_resp, 
  output        io_deq_bits_last 
);
  reg [63:0] _T_data [0:1]; 
  reg [63:0] _RAND_0;
  wire [63:0] _T_data__T_18_data; 
  wire  _T_data__T_18_addr; 
  wire [63:0] _T_data__T_10_data; 
  wire  _T_data__T_10_addr; 
  wire  _T_data__T_10_mask; 
  wire  _T_data__T_10_en; 
  reg [1:0] _T_resp [0:1]; 
  reg [31:0] _RAND_1;
  wire [1:0] _T_resp__T_18_data; 
  wire  _T_resp__T_18_addr; 
  wire [1:0] _T_resp__T_10_data; 
  wire  _T_resp__T_10_addr; 
  wire  _T_resp__T_10_mask; 
  wire  _T_resp__T_10_en; 
  reg  _T_last [0:1]; 
  reg [31:0] _RAND_2;
  wire  _T_last__T_18_data; 
  wire  _T_last__T_18_addr; 
  wire  _T_last__T_10_data; 
  wire  _T_last__T_10_addr; 
  wire  _T_last__T_10_mask; 
  wire  _T_last__T_10_en; 
  reg  value; 
  reg [31:0] _RAND_3;
  reg  value_1; 
  reg [31:0] _RAND_4;
  reg  _T_1; 
  reg [31:0] _RAND_5;
  wire  _T_2; 
  wire  _T_3; 
  wire  _T_4; 
  wire  _T_5; 
  wire  _T_6; 
  wire  _T_8; 
  wire  _T_12; 
  wire  _T_14; 
  wire  _T_15; 
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; 
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_resp__T_18_addr = value_1;
  assign _T_resp__T_18_data = _T_resp[_T_resp__T_18_addr]; 
  assign _T_resp__T_10_data = io_enq_bits_resp;
  assign _T_resp__T_10_addr = value;
  assign _T_resp__T_10_mask = 1'h1;
  assign _T_resp__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; 
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; 
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_4 = _T_2 & _T_3; 
  assign _T_5 = _T_2 & _T_1; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _T_12 = value + 1'h1; 
  assign _T_14 = value_1 + 1'h1; 
  assign _T_15 = _T_6 != _T_8; 
  assign io_enq_ready = _T_5 == 1'h0; 
  assign io_deq_valid = _T_4 == 1'h0; 
  assign io_deq_bits_data = _T_data__T_18_data; 
  assign io_deq_bits_resp = _T_resp__T_18_data; 
  assign io_deq_bits_last = _T_last__T_18_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_resp[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; 
    end
    if(_T_resp__T_10_en & _T_resp__T_10_mask) begin
      _T_resp[_T_resp__T_10_addr] <= _T_resp__T_10_data; 
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; 
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (_T_6) begin
        value <= _T_12;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (_T_8) begin
        value_1 <= _T_14;
      end
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_15) begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module dual_Queue_53( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [15:0] io_enq_bits, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [15:0] io_deq_bits 
);
  reg [15:0] _T [0:127]; 
  reg [31:0] _RAND_0;
  wire [15:0] _T__T_18_data; 
  wire [6:0] _T__T_18_addr; 
  wire [15:0] _T__T_10_data; 
  wire [6:0] _T__T_10_addr; 
  wire  _T__T_10_mask; 
  wire  _T__T_10_en; 
  reg [6:0] value; 
  reg [31:0] _RAND_1;
  reg [6:0] value_1; 
  reg [31:0] _RAND_2;
  reg  _T_1; 
  reg [31:0] _RAND_3;
  wire  _T_2; 
  wire  _T_3; 
  wire  _T_4; 
  wire  _T_5; 
  wire  _T_6; 
  wire  _T_8; 
  wire [6:0] _T_12; 
  wire [6:0] _T_14; 
  wire  _T_15; 
  assign _T__T_18_addr = value_1;
  assign _T__T_18_data = _T[_T__T_18_addr]; 
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = value;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; 
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_4 = _T_2 & _T_3; 
  assign _T_5 = _T_2 & _T_1; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _T_12 = value + 7'h1; 
  assign _T_14 = value_1 + 7'h1; 
  assign _T_15 = _T_6 != _T_8; 
  assign io_enq_ready = _T_5 == 1'h0; 
  assign io_deq_valid = _T_4 == 1'h0; 
  assign io_deq_bits = _T__T_18_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    _T[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; 
    end
    if (reset) begin
      value <= 7'h0;
    end else begin
      if (_T_6) begin
        value <= _T_12;
      end
    end
    if (reset) begin
      value_1 <= 7'h0;
    end else begin
      if (_T_8) begin
        value_1 <= _T_14;
      end
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_15) begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module dual_Queue_55( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [63:0] io_enq_bits_data, 
  input  [1:0]  io_enq_bits_resp, 
  input  [15:0] io_enq_bits_user, 
  input         io_enq_bits_last, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [63:0] io_deq_bits_data, 
  output [1:0]  io_deq_bits_resp, 
  output [15:0] io_deq_bits_user, 
  output        io_deq_bits_last 
);
  reg [63:0] _T_data [0:7]; 
  reg [63:0] _RAND_0;
  wire [63:0] _T_data__T_18_data; 
  wire [2:0] _T_data__T_18_addr; 
  wire [63:0] _T_data__T_10_data; 
  wire [2:0] _T_data__T_10_addr; 
  wire  _T_data__T_10_mask; 
  wire  _T_data__T_10_en; 
  reg [1:0] _T_resp [0:7]; 
  reg [31:0] _RAND_1;
  wire [1:0] _T_resp__T_18_data; 
  wire [2:0] _T_resp__T_18_addr; 
  wire [1:0] _T_resp__T_10_data; 
  wire [2:0] _T_resp__T_10_addr; 
  wire  _T_resp__T_10_mask; 
  wire  _T_resp__T_10_en; 
  reg [15:0] _T_user [0:7]; 
  reg [31:0] _RAND_2;
  wire [15:0] _T_user__T_18_data; 
  wire [2:0] _T_user__T_18_addr; 
  wire [15:0] _T_user__T_10_data; 
  wire [2:0] _T_user__T_10_addr; 
  wire  _T_user__T_10_mask; 
  wire  _T_user__T_10_en; 
  reg  _T_last [0:7]; 
  reg [31:0] _RAND_3;
  wire  _T_last__T_18_data; 
  wire [2:0] _T_last__T_18_addr; 
  wire  _T_last__T_10_data; 
  wire [2:0] _T_last__T_10_addr; 
  wire  _T_last__T_10_mask; 
  wire  _T_last__T_10_en; 
  reg [2:0] value; 
  reg [31:0] _RAND_4;
  reg [2:0] value_1; 
  reg [31:0] _RAND_5;
  reg  _T_1; 
  reg [31:0] _RAND_6;
  wire  _T_2; 
  wire  _T_3; 
  wire  _T_4; 
  wire  _T_5; 
  wire  _T_6; 
  wire  _T_8; 
  wire [2:0] _T_12; 
  wire [2:0] _T_14; 
  wire  _T_15; 
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; 
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_resp__T_18_addr = value_1;
  assign _T_resp__T_18_data = _T_resp[_T_resp__T_18_addr]; 
  assign _T_resp__T_10_data = io_enq_bits_resp;
  assign _T_resp__T_10_addr = value;
  assign _T_resp__T_10_mask = 1'h1;
  assign _T_resp__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_user__T_18_addr = value_1;
  assign _T_user__T_18_data = _T_user[_T_user__T_18_addr]; 
  assign _T_user__T_10_data = io_enq_bits_user;
  assign _T_user__T_10_addr = value;
  assign _T_user__T_10_mask = 1'h1;
  assign _T_user__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; 
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; 
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_4 = _T_2 & _T_3; 
  assign _T_5 = _T_2 & _T_1; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _T_12 = value + 3'h1; 
  assign _T_14 = value_1 + 3'h1; 
  assign _T_15 = _T_6 != _T_8; 
  assign io_enq_ready = _T_5 == 1'h0; 
  assign io_deq_valid = _T_4 == 1'h0; 
  assign io_deq_bits_data = _T_data__T_18_data; 
  assign io_deq_bits_resp = _T_resp__T_18_data; 
  assign io_deq_bits_user = _T_user__T_18_data; 
  assign io_deq_bits_last = _T_last__T_18_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    _T_resp[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    _T_user[initvar] = _RAND_2[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    _T_last[initvar] = _RAND_3[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value_1 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; 
    end
    if(_T_resp__T_10_en & _T_resp__T_10_mask) begin
      _T_resp[_T_resp__T_10_addr] <= _T_resp__T_10_data; 
    end
    if(_T_user__T_10_en & _T_user__T_10_mask) begin
      _T_user[_T_user__T_10_addr] <= _T_user__T_10_data; 
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; 
    end
    if (reset) begin
      value <= 3'h0;
    end else begin
      if (_T_6) begin
        value <= _T_12;
      end
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else begin
      if (_T_8) begin
        value_1 <= _T_14;
      end
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_15) begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module dual_Queue_57( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [4:0]  io_enq_bits_id, 
  input  [30:0] io_enq_bits_addr, 
  input  [7:0]  io_enq_bits_len, 
  input  [2:0]  io_enq_bits_size, 
  input  [10:0] io_enq_bits_user, 
  input         io_enq_bits_wen, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [4:0]  io_deq_bits_id, 
  output [30:0] io_deq_bits_addr, 
  output [7:0]  io_deq_bits_len, 
  output [2:0]  io_deq_bits_size, 
  output [1:0]  io_deq_bits_burst, 
  output        io_deq_bits_lock, 
  output [3:0]  io_deq_bits_cache, 
  output [2:0]  io_deq_bits_prot, 
  output [3:0]  io_deq_bits_qos, 
  output [10:0] io_deq_bits_user, 
  output [63:0] io_deq_bits_instret, 
  output        io_deq_bits_wen 
);
  reg [4:0] _T_id [0:0]; 
  reg [31:0] _RAND_0;
  wire [4:0] _T_id__T_14_data; 
  wire  _T_id__T_14_addr; 
  wire [4:0] _T_id__T_10_data; 
  wire  _T_id__T_10_addr; 
  wire  _T_id__T_10_mask; 
  wire  _T_id__T_10_en; 
  reg [30:0] _T_addr [0:0]; 
  reg [31:0] _RAND_1;
  wire [30:0] _T_addr__T_14_data; 
  wire  _T_addr__T_14_addr; 
  wire [30:0] _T_addr__T_10_data; 
  wire  _T_addr__T_10_addr; 
  wire  _T_addr__T_10_mask; 
  wire  _T_addr__T_10_en; 
  reg [7:0] _T_len [0:0]; 
  reg [31:0] _RAND_2;
  wire [7:0] _T_len__T_14_data; 
  wire  _T_len__T_14_addr; 
  wire [7:0] _T_len__T_10_data; 
  wire  _T_len__T_10_addr; 
  wire  _T_len__T_10_mask; 
  wire  _T_len__T_10_en; 
  reg [2:0] _T_size [0:0]; 
  reg [31:0] _RAND_3;
  wire [2:0] _T_size__T_14_data; 
  wire  _T_size__T_14_addr; 
  wire [2:0] _T_size__T_10_data; 
  wire  _T_size__T_10_addr; 
  wire  _T_size__T_10_mask; 
  wire  _T_size__T_10_en; 
  reg [1:0] _T_burst [0:0]; 
  reg [31:0] _RAND_4;
  wire [1:0] _T_burst__T_14_data; 
  wire  _T_burst__T_14_addr; 
  wire [1:0] _T_burst__T_10_data; 
  wire  _T_burst__T_10_addr; 
  wire  _T_burst__T_10_mask; 
  wire  _T_burst__T_10_en; 
  reg  _T_lock [0:0]; 
  reg [31:0] _RAND_5;
  wire  _T_lock__T_14_data; 
  wire  _T_lock__T_14_addr; 
  wire  _T_lock__T_10_data; 
  wire  _T_lock__T_10_addr; 
  wire  _T_lock__T_10_mask; 
  wire  _T_lock__T_10_en; 
  reg [3:0] _T_cache [0:0]; 
  reg [31:0] _RAND_6;
  wire [3:0] _T_cache__T_14_data; 
  wire  _T_cache__T_14_addr; 
  wire [3:0] _T_cache__T_10_data; 
  wire  _T_cache__T_10_addr; 
  wire  _T_cache__T_10_mask; 
  wire  _T_cache__T_10_en; 
  reg [2:0] _T_prot [0:0]; 
  reg [31:0] _RAND_7;
  wire [2:0] _T_prot__T_14_data; 
  wire  _T_prot__T_14_addr; 
  wire [2:0] _T_prot__T_10_data; 
  wire  _T_prot__T_10_addr; 
  wire  _T_prot__T_10_mask; 
  wire  _T_prot__T_10_en; 
  reg [3:0] _T_qos [0:0]; 
  reg [31:0] _RAND_8;
  wire [3:0] _T_qos__T_14_data; 
  wire  _T_qos__T_14_addr; 
  wire [3:0] _T_qos__T_10_data; 
  wire  _T_qos__T_10_addr; 
  wire  _T_qos__T_10_mask; 
  wire  _T_qos__T_10_en; 
  reg [10:0] _T_user [0:0]; 
  reg [31:0] _RAND_9;
  wire [10:0] _T_user__T_14_data; 
  wire  _T_user__T_14_addr; 
  wire [10:0] _T_user__T_10_data; 
  wire  _T_user__T_10_addr; 
  wire  _T_user__T_10_mask; 
  wire  _T_user__T_10_en; 
  reg [63:0] _T_instret [0:0]; 
  reg [63:0] _RAND_10;
  wire [63:0] _T_instret__T_14_data; 
  wire  _T_instret__T_14_addr; 
  wire [63:0] _T_instret__T_10_data; 
  wire  _T_instret__T_10_addr; 
  wire  _T_instret__T_10_mask; 
  wire  _T_instret__T_10_en; 
  reg  _T_wen [0:0]; 
  reg [31:0] _RAND_11;
  wire  _T_wen__T_14_data; 
  wire  _T_wen__T_14_addr; 
  wire  _T_wen__T_10_data; 
  wire  _T_wen__T_10_addr; 
  wire  _T_wen__T_10_mask; 
  wire  _T_wen__T_10_en; 
  reg  _T_1; 
  reg [31:0] _RAND_12;
  wire  _T_3; 
  wire  _T_6; 
  wire  _T_8; 
  wire  _GEN_18; 
  wire  _GEN_32; 
  wire  _GEN_31; 
  wire  _T_11; 
  wire  _T_12; 
  assign _T_id__T_14_addr = 1'h0;
  assign _T_id__T_14_data = _T_id[_T_id__T_14_addr]; 
  assign _T_id__T_10_data = io_enq_bits_id;
  assign _T_id__T_10_addr = 1'h0;
  assign _T_id__T_10_mask = 1'h1;
  assign _T_id__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_addr__T_14_addr = 1'h0;
  assign _T_addr__T_14_data = _T_addr[_T_addr__T_14_addr]; 
  assign _T_addr__T_10_data = io_enq_bits_addr;
  assign _T_addr__T_10_addr = 1'h0;
  assign _T_addr__T_10_mask = 1'h1;
  assign _T_addr__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_len__T_14_addr = 1'h0;
  assign _T_len__T_14_data = _T_len[_T_len__T_14_addr]; 
  assign _T_len__T_10_data = io_enq_bits_len;
  assign _T_len__T_10_addr = 1'h0;
  assign _T_len__T_10_mask = 1'h1;
  assign _T_len__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_size__T_14_addr = 1'h0;
  assign _T_size__T_14_data = _T_size[_T_size__T_14_addr]; 
  assign _T_size__T_10_data = io_enq_bits_size;
  assign _T_size__T_10_addr = 1'h0;
  assign _T_size__T_10_mask = 1'h1;
  assign _T_size__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_burst__T_14_addr = 1'h0;
  assign _T_burst__T_14_data = _T_burst[_T_burst__T_14_addr]; 
  assign _T_burst__T_10_data = 2'h1;
  assign _T_burst__T_10_addr = 1'h0;
  assign _T_burst__T_10_mask = 1'h1;
  assign _T_burst__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_lock__T_14_addr = 1'h0;
  assign _T_lock__T_14_data = _T_lock[_T_lock__T_14_addr]; 
  assign _T_lock__T_10_data = 1'h0;
  assign _T_lock__T_10_addr = 1'h0;
  assign _T_lock__T_10_mask = 1'h1;
  assign _T_lock__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_cache__T_14_addr = 1'h0;
  assign _T_cache__T_14_data = _T_cache[_T_cache__T_14_addr]; 
  assign _T_cache__T_10_data = 4'h0;
  assign _T_cache__T_10_addr = 1'h0;
  assign _T_cache__T_10_mask = 1'h1;
  assign _T_cache__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_prot__T_14_addr = 1'h0;
  assign _T_prot__T_14_data = _T_prot[_T_prot__T_14_addr]; 
  assign _T_prot__T_10_data = 3'h1;
  assign _T_prot__T_10_addr = 1'h0;
  assign _T_prot__T_10_mask = 1'h1;
  assign _T_prot__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_qos__T_14_addr = 1'h0;
  assign _T_qos__T_14_data = _T_qos[_T_qos__T_14_addr]; 
  assign _T_qos__T_10_data = 4'h0;
  assign _T_qos__T_10_addr = 1'h0;
  assign _T_qos__T_10_mask = 1'h1;
  assign _T_qos__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_user__T_14_addr = 1'h0;
  assign _T_user__T_14_data = _T_user[_T_user__T_14_addr]; 
  assign _T_user__T_10_data = io_enq_bits_user;
  assign _T_user__T_10_addr = 1'h0;
  assign _T_user__T_10_mask = 1'h1;
  assign _T_user__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_instret__T_14_addr = 1'h0;
  assign _T_instret__T_14_data = _T_instret[_T_instret__T_14_addr]; 
  assign _T_instret__T_10_data = 64'h0;
  assign _T_instret__T_10_addr = 1'h0;
  assign _T_instret__T_10_mask = 1'h1;
  assign _T_instret__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_wen__T_14_addr = 1'h0;
  assign _T_wen__T_14_data = _T_wen[_T_wen__T_14_addr]; 
  assign _T_wen__T_10_data = io_enq_bits_wen;
  assign _T_wen__T_10_addr = 1'h0;
  assign _T_wen__T_10_mask = 1'h1;
  assign _T_wen__T_10_en = _T_3 ? _GEN_18 : _T_6;
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _GEN_18 = io_deq_ready ? 1'h0 : _T_6; 
  assign _GEN_32 = _T_3 ? _GEN_18 : _T_6; 
  assign _GEN_31 = _T_3 ? 1'h0 : _T_8; 
  assign _T_11 = _GEN_32 != _GEN_31; 
  assign _T_12 = _T_3 == 1'h0; 
  assign io_enq_ready = _T_1 == 1'h0; 
  assign io_deq_valid = io_enq_valid ? 1'h1 : _T_12; 
  assign io_deq_bits_id = _T_3 ? io_enq_bits_id : _T_id__T_14_data; 
  assign io_deq_bits_addr = _T_3 ? io_enq_bits_addr : _T_addr__T_14_data; 
  assign io_deq_bits_len = _T_3 ? io_enq_bits_len : _T_len__T_14_data; 
  assign io_deq_bits_size = _T_3 ? io_enq_bits_size : _T_size__T_14_data; 
  assign io_deq_bits_burst = _T_3 ? 2'h1 : _T_burst__T_14_data; 
  assign io_deq_bits_lock = _T_3 ? 1'h0 : _T_lock__T_14_data; 
  assign io_deq_bits_cache = _T_3 ? 4'h0 : _T_cache__T_14_data; 
  assign io_deq_bits_prot = _T_3 ? 3'h1 : _T_prot__T_14_data; 
  assign io_deq_bits_qos = _T_3 ? 4'h0 : _T_qos__T_14_data; 
  assign io_deq_bits_user = _T_3 ? io_enq_bits_user : _T_user__T_14_data; 
  assign io_deq_bits_instret = _T_3 ? 64'h0 : _T_instret__T_14_data; 
  assign io_deq_bits_wen = _T_3 ? io_enq_bits_wen : _T_wen__T_14_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_id[initvar] = _RAND_0[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_addr[initvar] = _RAND_1[30:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_len[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_size[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_burst[initvar] = _RAND_4[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_lock[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_cache[initvar] = _RAND_6[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_prot[initvar] = _RAND_7[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_qos[initvar] = _RAND_8[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_user[initvar] = _RAND_9[10:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_10 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_instret[initvar] = _RAND_10[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_11 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_wen[initvar] = _RAND_11[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_1 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T_id__T_10_en & _T_id__T_10_mask) begin
      _T_id[_T_id__T_10_addr] <= _T_id__T_10_data; 
    end
    if(_T_addr__T_10_en & _T_addr__T_10_mask) begin
      _T_addr[_T_addr__T_10_addr] <= _T_addr__T_10_data; 
    end
    if(_T_len__T_10_en & _T_len__T_10_mask) begin
      _T_len[_T_len__T_10_addr] <= _T_len__T_10_data; 
    end
    if(_T_size__T_10_en & _T_size__T_10_mask) begin
      _T_size[_T_size__T_10_addr] <= _T_size__T_10_data; 
    end
    if(_T_burst__T_10_en & _T_burst__T_10_mask) begin
      _T_burst[_T_burst__T_10_addr] <= _T_burst__T_10_data; 
    end
    if(_T_lock__T_10_en & _T_lock__T_10_mask) begin
      _T_lock[_T_lock__T_10_addr] <= _T_lock__T_10_data; 
    end
    if(_T_cache__T_10_en & _T_cache__T_10_mask) begin
      _T_cache[_T_cache__T_10_addr] <= _T_cache__T_10_data; 
    end
    if(_T_prot__T_10_en & _T_prot__T_10_mask) begin
      _T_prot[_T_prot__T_10_addr] <= _T_prot__T_10_data; 
    end
    if(_T_qos__T_10_en & _T_qos__T_10_mask) begin
      _T_qos[_T_qos__T_10_addr] <= _T_qos__T_10_data; 
    end
    if(_T_user__T_10_en & _T_user__T_10_mask) begin
      _T_user[_T_user__T_10_addr] <= _T_user__T_10_data; 
    end
    if(_T_instret__T_10_en & _T_instret__T_10_mask) begin
      _T_instret[_T_instret__T_10_addr] <= _T_instret__T_10_data; 
    end
    if(_T_wen__T_10_en & _T_wen__T_10_mask) begin
      _T_wen[_T_wen__T_10_addr] <= _T_wen__T_10_data; 
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_3) begin
          if (io_deq_ready) begin
            _T_1 <= 1'h0;
          end else begin
            _T_1 <= _T_6;
          end
        end else begin
          _T_1 <= _T_6;
        end
      end
    end
  end
endmodule
module dual_Queue_58( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input         io_enq_bits_id, 
  input  [63:0] io_enq_bits_data, 
  input  [1:0]  io_enq_bits_resp, 
  input         io_enq_bits_last, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output        io_deq_bits_id, 
  output [63:0] io_deq_bits_data, 
  output [1:0]  io_deq_bits_resp, 
  output        io_deq_bits_last 
);
  reg  _T_id [0:0]; 
  reg [31:0] _RAND_0;
  wire  _T_id__T_14_data; 
  wire  _T_id__T_14_addr; 
  wire  _T_id__T_10_data; 
  wire  _T_id__T_10_addr; 
  wire  _T_id__T_10_mask; 
  wire  _T_id__T_10_en; 
  reg [63:0] _T_data [0:0]; 
  reg [63:0] _RAND_1;
  wire [63:0] _T_data__T_14_data; 
  wire  _T_data__T_14_addr; 
  wire [63:0] _T_data__T_10_data; 
  wire  _T_data__T_10_addr; 
  wire  _T_data__T_10_mask; 
  wire  _T_data__T_10_en; 
  reg [1:0] _T_resp [0:0]; 
  reg [31:0] _RAND_2;
  wire [1:0] _T_resp__T_14_data; 
  wire  _T_resp__T_14_addr; 
  wire [1:0] _T_resp__T_10_data; 
  wire  _T_resp__T_10_addr; 
  wire  _T_resp__T_10_mask; 
  wire  _T_resp__T_10_en; 
  reg  _T_last [0:0]; 
  reg [31:0] _RAND_3;
  wire  _T_last__T_14_data; 
  wire  _T_last__T_14_addr; 
  wire  _T_last__T_10_data; 
  wire  _T_last__T_10_addr; 
  wire  _T_last__T_10_mask; 
  wire  _T_last__T_10_en; 
  reg  _T_1; 
  reg [31:0] _RAND_4;
  wire  _T_3; 
  wire  _T_6; 
  wire  _T_8; 
  wire  _GEN_10; 
  wire  _GEN_16; 
  wire  _GEN_15; 
  wire  _T_11; 
  wire  _T_12; 
  assign _T_id__T_14_addr = 1'h0;
  assign _T_id__T_14_data = _T_id[_T_id__T_14_addr]; 
  assign _T_id__T_10_data = io_enq_bits_id;
  assign _T_id__T_10_addr = 1'h0;
  assign _T_id__T_10_mask = 1'h1;
  assign _T_id__T_10_en = _T_3 ? _GEN_10 : _T_6;
  assign _T_data__T_14_addr = 1'h0;
  assign _T_data__T_14_data = _T_data[_T_data__T_14_addr]; 
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = 1'h0;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = _T_3 ? _GEN_10 : _T_6;
  assign _T_resp__T_14_addr = 1'h0;
  assign _T_resp__T_14_data = _T_resp[_T_resp__T_14_addr]; 
  assign _T_resp__T_10_data = io_enq_bits_resp;
  assign _T_resp__T_10_addr = 1'h0;
  assign _T_resp__T_10_mask = 1'h1;
  assign _T_resp__T_10_en = _T_3 ? _GEN_10 : _T_6;
  assign _T_last__T_14_addr = 1'h0;
  assign _T_last__T_14_data = _T_last[_T_last__T_14_addr]; 
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = 1'h0;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = _T_3 ? _GEN_10 : _T_6;
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _GEN_10 = io_deq_ready ? 1'h0 : _T_6; 
  assign _GEN_16 = _T_3 ? _GEN_10 : _T_6; 
  assign _GEN_15 = _T_3 ? 1'h0 : _T_8; 
  assign _T_11 = _GEN_16 != _GEN_15; 
  assign _T_12 = _T_3 == 1'h0; 
  assign io_enq_ready = _T_1 == 1'h0; 
  assign io_deq_valid = io_enq_valid ? 1'h1 : _T_12; 
  assign io_deq_bits_id = _T_3 ? io_enq_bits_id : _T_id__T_14_data; 
  assign io_deq_bits_data = _T_3 ? io_enq_bits_data : _T_data__T_14_data; 
  assign io_deq_bits_resp = _T_3 ? io_enq_bits_resp : _T_resp__T_14_data; 
  assign io_deq_bits_last = _T_3 ? io_enq_bits_last : _T_last__T_14_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_id[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_data[initvar] = _RAND_1[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_resp[initvar] = _RAND_2[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_last[initvar] = _RAND_3[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T_id__T_10_en & _T_id__T_10_mask) begin
      _T_id[_T_id__T_10_addr] <= _T_id__T_10_data; 
    end
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; 
    end
    if(_T_resp__T_10_en & _T_resp__T_10_mask) begin
      _T_resp[_T_resp__T_10_addr] <= _T_resp__T_10_data; 
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; 
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_3) begin
          if (io_deq_ready) begin
            _T_1 <= 1'h0;
          end else begin
            _T_1 <= _T_6;
          end
        end else begin
          _T_1 <= _T_6;
        end
      end
    end
  end
endmodule
module dual_Queue_59( 
  input        clock, 
  input        reset, 
  output       io_enq_ready, 
  input        io_enq_valid, 
  input        io_enq_bits_id, 
  input  [1:0] io_enq_bits_resp, 
  input        io_deq_ready, 
  output       io_deq_valid, 
  output       io_deq_bits_id, 
  output [1:0] io_deq_bits_resp 
);
  reg  _T_id [0:0]; 
  reg [31:0] _RAND_0;
  wire  _T_id__T_14_data; 
  wire  _T_id__T_14_addr; 
  wire  _T_id__T_10_data; 
  wire  _T_id__T_10_addr; 
  wire  _T_id__T_10_mask; 
  wire  _T_id__T_10_en; 
  reg [1:0] _T_resp [0:0]; 
  reg [31:0] _RAND_1;
  wire [1:0] _T_resp__T_14_data; 
  wire  _T_resp__T_14_addr; 
  wire [1:0] _T_resp__T_10_data; 
  wire  _T_resp__T_10_addr; 
  wire  _T_resp__T_10_mask; 
  wire  _T_resp__T_10_en; 
  reg  _T_1; 
  reg [31:0] _RAND_2;
  wire  _T_3; 
  wire  _T_6; 
  wire  _T_8; 
  wire  _GEN_8; 
  wire  _GEN_12; 
  wire  _GEN_11; 
  wire  _T_11; 
  wire  _T_12; 
  assign _T_id__T_14_addr = 1'h0;
  assign _T_id__T_14_data = _T_id[_T_id__T_14_addr]; 
  assign _T_id__T_10_data = io_enq_bits_id;
  assign _T_id__T_10_addr = 1'h0;
  assign _T_id__T_10_mask = 1'h1;
  assign _T_id__T_10_en = _T_3 ? _GEN_8 : _T_6;
  assign _T_resp__T_14_addr = 1'h0;
  assign _T_resp__T_14_data = _T_resp[_T_resp__T_14_addr]; 
  assign _T_resp__T_10_data = io_enq_bits_resp;
  assign _T_resp__T_10_addr = 1'h0;
  assign _T_resp__T_10_mask = 1'h1;
  assign _T_resp__T_10_en = _T_3 ? _GEN_8 : _T_6;
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _GEN_8 = io_deq_ready ? 1'h0 : _T_6; 
  assign _GEN_12 = _T_3 ? _GEN_8 : _T_6; 
  assign _GEN_11 = _T_3 ? 1'h0 : _T_8; 
  assign _T_11 = _GEN_12 != _GEN_11; 
  assign _T_12 = _T_3 == 1'h0; 
  assign io_enq_ready = _T_1 == 1'h0; 
  assign io_deq_valid = io_enq_valid ? 1'h1 : _T_12; 
  assign io_deq_bits_id = _T_3 ? io_enq_bits_id : _T_id__T_14_data; 
  assign io_deq_bits_resp = _T_3 ? io_enq_bits_resp : _T_resp__T_14_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_id[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_resp[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T_id__T_10_en & _T_id__T_10_mask) begin
      _T_id[_T_id__T_10_addr] <= _T_id__T_10_data; 
    end
    if(_T_resp__T_10_en & _T_resp__T_10_mask) begin
      _T_resp[_T_resp__T_10_addr] <= _T_resp__T_10_data; 
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_3) begin
          if (io_deq_ready) begin
            _T_1 <= 1'h0;
          end else begin
            _T_1 <= _T_6;
          end
        end else begin
          _T_1 <= _T_6;
        end
      end
    end
  end
endmodule
module dual_Queue_5( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [2:0]  io_enq_bits_opcode, 
  input  [2:0]  io_enq_bits_param, 
  input  [2:0]  io_enq_bits_size, 
  input  [2:0]  io_enq_bits_source, 
  input  [31:0] io_enq_bits_address, 
  input  [3:0]  io_enq_bits_mask, 
  input  [31:0] io_enq_bits_data, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [2:0]  io_deq_bits_opcode, 
  output [2:0]  io_deq_bits_param, 
  output [2:0]  io_deq_bits_size, 
  output [2:0]  io_deq_bits_source, 
  output [31:0] io_deq_bits_address, 
  output [3:0]  io_deq_bits_mask, 
  output [31:0] io_deq_bits_data 
);
  reg [2:0] _T_opcode [0:0]; 
  reg [31:0] _RAND_0;
  wire [2:0] _T_opcode__T_14_data; 
  wire  _T_opcode__T_14_addr; 
  wire [2:0] _T_opcode__T_10_data; 
  wire  _T_opcode__T_10_addr; 
  wire  _T_opcode__T_10_mask; 
  wire  _T_opcode__T_10_en; 
  reg [2:0] _T_param [0:0]; 
  reg [31:0] _RAND_1;
  wire [2:0] _T_param__T_14_data; 
  wire  _T_param__T_14_addr; 
  wire [2:0] _T_param__T_10_data; 
  wire  _T_param__T_10_addr; 
  wire  _T_param__T_10_mask; 
  wire  _T_param__T_10_en; 
  reg [2:0] _T_size [0:0]; 
  reg [31:0] _RAND_2;
  wire [2:0] _T_size__T_14_data; 
  wire  _T_size__T_14_addr; 
  wire [2:0] _T_size__T_10_data; 
  wire  _T_size__T_10_addr; 
  wire  _T_size__T_10_mask; 
  wire  _T_size__T_10_en; 
  reg [2:0] _T_source [0:0]; 
  reg [31:0] _RAND_3;
  wire [2:0] _T_source__T_14_data; 
  wire  _T_source__T_14_addr; 
  wire [2:0] _T_source__T_10_data; 
  wire  _T_source__T_10_addr; 
  wire  _T_source__T_10_mask; 
  wire  _T_source__T_10_en; 
  reg [31:0] _T_address [0:0]; 
  reg [31:0] _RAND_4;
  wire [31:0] _T_address__T_14_data; 
  wire  _T_address__T_14_addr; 
  wire [31:0] _T_address__T_10_data; 
  wire  _T_address__T_10_addr; 
  wire  _T_address__T_10_mask; 
  wire  _T_address__T_10_en; 
  reg [3:0] _T_mask [0:0]; 
  reg [31:0] _RAND_5;
  wire [3:0] _T_mask__T_14_data; 
  wire  _T_mask__T_14_addr; 
  wire [3:0] _T_mask__T_10_data; 
  wire  _T_mask__T_10_addr; 
  wire  _T_mask__T_10_mask; 
  wire  _T_mask__T_10_en; 
  reg [31:0] _T_data [0:0]; 
  reg [31:0] _RAND_6;
  wire [31:0] _T_data__T_14_data; 
  wire  _T_data__T_14_addr; 
  wire [31:0] _T_data__T_10_data; 
  wire  _T_data__T_10_addr; 
  wire  _T_data__T_10_mask; 
  wire  _T_data__T_10_en; 
  reg  _T_1; 
  reg [31:0] _RAND_7;
  wire  _T_3; 
  wire  _T_6; 
  wire  _T_8; 
  wire  _GEN_16; 
  wire  _GEN_28; 
  wire  _GEN_27; 
  wire  _T_11; 
  wire  _T_12; 
  assign _T_opcode__T_14_addr = 1'h0;
  assign _T_opcode__T_14_data = _T_opcode[_T_opcode__T_14_addr]; 
  assign _T_opcode__T_10_data = io_enq_bits_opcode;
  assign _T_opcode__T_10_addr = 1'h0;
  assign _T_opcode__T_10_mask = 1'h1;
  assign _T_opcode__T_10_en = _T_3 ? _GEN_16 : _T_6;
  assign _T_param__T_14_addr = 1'h0;
  assign _T_param__T_14_data = _T_param[_T_param__T_14_addr]; 
  assign _T_param__T_10_data = io_enq_bits_param;
  assign _T_param__T_10_addr = 1'h0;
  assign _T_param__T_10_mask = 1'h1;
  assign _T_param__T_10_en = _T_3 ? _GEN_16 : _T_6;
  assign _T_size__T_14_addr = 1'h0;
  assign _T_size__T_14_data = _T_size[_T_size__T_14_addr]; 
  assign _T_size__T_10_data = io_enq_bits_size;
  assign _T_size__T_10_addr = 1'h0;
  assign _T_size__T_10_mask = 1'h1;
  assign _T_size__T_10_en = _T_3 ? _GEN_16 : _T_6;
  assign _T_source__T_14_addr = 1'h0;
  assign _T_source__T_14_data = _T_source[_T_source__T_14_addr]; 
  assign _T_source__T_10_data = io_enq_bits_source;
  assign _T_source__T_10_addr = 1'h0;
  assign _T_source__T_10_mask = 1'h1;
  assign _T_source__T_10_en = _T_3 ? _GEN_16 : _T_6;
  assign _T_address__T_14_addr = 1'h0;
  assign _T_address__T_14_data = _T_address[_T_address__T_14_addr]; 
  assign _T_address__T_10_data = io_enq_bits_address;
  assign _T_address__T_10_addr = 1'h0;
  assign _T_address__T_10_mask = 1'h1;
  assign _T_address__T_10_en = _T_3 ? _GEN_16 : _T_6;
  assign _T_mask__T_14_addr = 1'h0;
  assign _T_mask__T_14_data = _T_mask[_T_mask__T_14_addr]; 
  assign _T_mask__T_10_data = io_enq_bits_mask;
  assign _T_mask__T_10_addr = 1'h0;
  assign _T_mask__T_10_mask = 1'h1;
  assign _T_mask__T_10_en = _T_3 ? _GEN_16 : _T_6;
  assign _T_data__T_14_addr = 1'h0;
  assign _T_data__T_14_data = _T_data[_T_data__T_14_addr]; 
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = 1'h0;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = _T_3 ? _GEN_16 : _T_6;
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _GEN_16 = io_deq_ready ? 1'h0 : _T_6; 
  assign _GEN_28 = _T_3 ? _GEN_16 : _T_6; 
  assign _GEN_27 = _T_3 ? 1'h0 : _T_8; 
  assign _T_11 = _GEN_28 != _GEN_27; 
  assign _T_12 = _T_3 == 1'h0; 
  assign io_enq_ready = _T_1 == 1'h0; 
  assign io_deq_valid = io_enq_valid ? 1'h1 : _T_12; 
  assign io_deq_bits_opcode = _T_3 ? io_enq_bits_opcode : _T_opcode__T_14_data; 
  assign io_deq_bits_param = _T_3 ? io_enq_bits_param : _T_param__T_14_data; 
  assign io_deq_bits_size = _T_3 ? io_enq_bits_size : _T_size__T_14_data; 
  assign io_deq_bits_source = _T_3 ? io_enq_bits_source : _T_source__T_14_data; 
  assign io_deq_bits_address = _T_3 ? io_enq_bits_address : _T_address__T_14_data; 
  assign io_deq_bits_mask = _T_3 ? io_enq_bits_mask : _T_mask__T_14_data; 
  assign io_deq_bits_data = _T_3 ? io_enq_bits_data : _T_data__T_14_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_param[initvar] = _RAND_1[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_size[initvar] = _RAND_2[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_source[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_address[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_mask[initvar] = _RAND_5[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_data[initvar] = _RAND_6[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_1 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T_opcode__T_10_en & _T_opcode__T_10_mask) begin
      _T_opcode[_T_opcode__T_10_addr] <= _T_opcode__T_10_data; 
    end
    if(_T_param__T_10_en & _T_param__T_10_mask) begin
      _T_param[_T_param__T_10_addr] <= _T_param__T_10_data; 
    end
    if(_T_size__T_10_en & _T_size__T_10_mask) begin
      _T_size[_T_size__T_10_addr] <= _T_size__T_10_data; 
    end
    if(_T_source__T_10_en & _T_source__T_10_mask) begin
      _T_source[_T_source__T_10_addr] <= _T_source__T_10_data; 
    end
    if(_T_address__T_10_en & _T_address__T_10_mask) begin
      _T_address[_T_address__T_10_addr] <= _T_address__T_10_data; 
    end
    if(_T_mask__T_10_en & _T_mask__T_10_mask) begin
      _T_mask[_T_mask__T_10_addr] <= _T_mask__T_10_data; 
    end
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; 
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_3) begin
          if (io_deq_ready) begin
            _T_1 <= 1'h0;
          end else begin
            _T_1 <= _T_6;
          end
        end else begin
          _T_1 <= _T_6;
        end
      end
    end
  end
endmodule
module dual_Queue_60( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [16:0] io_enq_bits, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [16:0] io_deq_bits 
);
  reg [16:0] _T [0:1]; 
  reg [31:0] _RAND_0;
  wire [16:0] _T__T_18_data; 
  wire  _T__T_18_addr; 
  wire [16:0] _T__T_10_data; 
  wire  _T__T_10_addr; 
  wire  _T__T_10_mask; 
  wire  _T__T_10_en; 
  reg  value; 
  reg [31:0] _RAND_1;
  reg  value_1; 
  reg [31:0] _RAND_2;
  reg  _T_1; 
  reg [31:0] _RAND_3;
  wire  _T_2; 
  wire  _T_3; 
  wire  _T_4; 
  wire  _T_5; 
  wire  _T_6; 
  wire  _T_8; 
  wire  _T_12; 
  wire  _T_14; 
  wire  _T_15; 
  assign _T__T_18_addr = value_1;
  assign _T__T_18_data = _T[_T__T_18_addr]; 
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = value;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; 
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_4 = _T_2 & _T_3; 
  assign _T_5 = _T_2 & _T_1; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _T_12 = value + 1'h1; 
  assign _T_14 = value_1 + 1'h1; 
  assign _T_15 = _T_6 != _T_8; 
  assign io_enq_ready = _T_5 == 1'h0; 
  assign io_deq_valid = _T_4 == 1'h0; 
  assign io_deq_bits = _T__T_18_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T[initvar] = _RAND_0[16:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; 
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (_T_6) begin
        value <= _T_12;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (_T_8) begin
        value_1 <= _T_14;
      end
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_15) begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module dual_Queue_64( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input         io_enq_bits_id, 
  input  [31:0] io_enq_bits_addr, 
  input  [7:0]  io_enq_bits_len, 
  input  [2:0]  io_enq_bits_size, 
  input  [1:0]  io_enq_bits_burst, 
  input  [15:0] io_enq_bits_user, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output        io_deq_bits_id, 
  output [31:0] io_deq_bits_addr, 
  output [7:0]  io_deq_bits_len, 
  output [2:0]  io_deq_bits_size, 
  output [1:0]  io_deq_bits_burst, 
  output [15:0] io_deq_bits_user 
);
  reg  _T_id [0:0]; 
  reg [31:0] _RAND_0;
  wire  _T_id__T_14_data; 
  wire  _T_id__T_14_addr; 
  wire  _T_id__T_10_data; 
  wire  _T_id__T_10_addr; 
  wire  _T_id__T_10_mask; 
  wire  _T_id__T_10_en; 
  reg [31:0] _T_addr [0:0]; 
  reg [31:0] _RAND_1;
  wire [31:0] _T_addr__T_14_data; 
  wire  _T_addr__T_14_addr; 
  wire [31:0] _T_addr__T_10_data; 
  wire  _T_addr__T_10_addr; 
  wire  _T_addr__T_10_mask; 
  wire  _T_addr__T_10_en; 
  reg [7:0] _T_len [0:0]; 
  reg [31:0] _RAND_2;
  wire [7:0] _T_len__T_14_data; 
  wire  _T_len__T_14_addr; 
  wire [7:0] _T_len__T_10_data; 
  wire  _T_len__T_10_addr; 
  wire  _T_len__T_10_mask; 
  wire  _T_len__T_10_en; 
  reg [2:0] _T_size [0:0]; 
  reg [31:0] _RAND_3;
  wire [2:0] _T_size__T_14_data; 
  wire  _T_size__T_14_addr; 
  wire [2:0] _T_size__T_10_data; 
  wire  _T_size__T_10_addr; 
  wire  _T_size__T_10_mask; 
  wire  _T_size__T_10_en; 
  reg [1:0] _T_burst [0:0]; 
  reg [31:0] _RAND_4;
  wire [1:0] _T_burst__T_14_data; 
  wire  _T_burst__T_14_addr; 
  wire [1:0] _T_burst__T_10_data; 
  wire  _T_burst__T_10_addr; 
  wire  _T_burst__T_10_mask; 
  wire  _T_burst__T_10_en; 
  reg [15:0] _T_user [0:0]; 
  reg [31:0] _RAND_5;
  wire [15:0] _T_user__T_14_data; 
  wire  _T_user__T_14_addr; 
  wire [15:0] _T_user__T_10_data; 
  wire  _T_user__T_10_addr; 
  wire  _T_user__T_10_mask; 
  wire  _T_user__T_10_en; 
  reg  _T_1; 
  reg [31:0] _RAND_6;
  wire  _T_3; 
  wire  _T_6; 
  wire  _T_8; 
  wire  _GEN_17; 
  wire  _GEN_30; 
  wire  _GEN_29; 
  wire  _T_11; 
  wire  _T_12; 
  assign _T_id__T_14_addr = 1'h0;
  assign _T_id__T_14_data = _T_id[_T_id__T_14_addr]; 
  assign _T_id__T_10_data = io_enq_bits_id;
  assign _T_id__T_10_addr = 1'h0;
  assign _T_id__T_10_mask = 1'h1;
  assign _T_id__T_10_en = _T_3 ? _GEN_17 : _T_6;
  assign _T_addr__T_14_addr = 1'h0;
  assign _T_addr__T_14_data = _T_addr[_T_addr__T_14_addr]; 
  assign _T_addr__T_10_data = io_enq_bits_addr;
  assign _T_addr__T_10_addr = 1'h0;
  assign _T_addr__T_10_mask = 1'h1;
  assign _T_addr__T_10_en = _T_3 ? _GEN_17 : _T_6;
  assign _T_len__T_14_addr = 1'h0;
  assign _T_len__T_14_data = _T_len[_T_len__T_14_addr]; 
  assign _T_len__T_10_data = io_enq_bits_len;
  assign _T_len__T_10_addr = 1'h0;
  assign _T_len__T_10_mask = 1'h1;
  assign _T_len__T_10_en = _T_3 ? _GEN_17 : _T_6;
  assign _T_size__T_14_addr = 1'h0;
  assign _T_size__T_14_data = _T_size[_T_size__T_14_addr]; 
  assign _T_size__T_10_data = io_enq_bits_size;
  assign _T_size__T_10_addr = 1'h0;
  assign _T_size__T_10_mask = 1'h1;
  assign _T_size__T_10_en = _T_3 ? _GEN_17 : _T_6;
  assign _T_burst__T_14_addr = 1'h0;
  assign _T_burst__T_14_data = _T_burst[_T_burst__T_14_addr]; 
  assign _T_burst__T_10_data = io_enq_bits_burst;
  assign _T_burst__T_10_addr = 1'h0;
  assign _T_burst__T_10_mask = 1'h1;
  assign _T_burst__T_10_en = _T_3 ? _GEN_17 : _T_6;
  assign _T_user__T_14_addr = 1'h0;
  assign _T_user__T_14_data = _T_user[_T_user__T_14_addr]; 
  assign _T_user__T_10_data = io_enq_bits_user;
  assign _T_user__T_10_addr = 1'h0;
  assign _T_user__T_10_mask = 1'h1;
  assign _T_user__T_10_en = _T_3 ? _GEN_17 : _T_6;
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _GEN_17 = io_deq_ready ? 1'h0 : _T_6; 
  assign _GEN_30 = _T_3 ? _GEN_17 : _T_6; 
  assign _GEN_29 = _T_3 ? 1'h0 : _T_8; 
  assign _T_11 = _GEN_30 != _GEN_29; 
  assign _T_12 = _T_3 == 1'h0; 
  assign io_enq_ready = _T_1 == 1'h0; 
  assign io_deq_valid = io_enq_valid ? 1'h1 : _T_12; 
  assign io_deq_bits_id = _T_3 ? io_enq_bits_id : _T_id__T_14_data; 
  assign io_deq_bits_addr = _T_3 ? io_enq_bits_addr : _T_addr__T_14_data; 
  assign io_deq_bits_len = _T_3 ? io_enq_bits_len : _T_len__T_14_data; 
  assign io_deq_bits_size = _T_3 ? io_enq_bits_size : _T_size__T_14_data; 
  assign io_deq_bits_burst = _T_3 ? io_enq_bits_burst : _T_burst__T_14_data; 
  assign io_deq_bits_user = _T_3 ? io_enq_bits_user : _T_user__T_14_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_id[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_addr[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_len[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_size[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_burst[initvar] = _RAND_4[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_user[initvar] = _RAND_5[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T_id__T_10_en & _T_id__T_10_mask) begin
      _T_id[_T_id__T_10_addr] <= _T_id__T_10_data; 
    end
    if(_T_addr__T_10_en & _T_addr__T_10_mask) begin
      _T_addr[_T_addr__T_10_addr] <= _T_addr__T_10_data; 
    end
    if(_T_len__T_10_en & _T_len__T_10_mask) begin
      _T_len[_T_len__T_10_addr] <= _T_len__T_10_data; 
    end
    if(_T_size__T_10_en & _T_size__T_10_mask) begin
      _T_size[_T_size__T_10_addr] <= _T_size__T_10_data; 
    end
    if(_T_burst__T_10_en & _T_burst__T_10_mask) begin
      _T_burst[_T_burst__T_10_addr] <= _T_burst__T_10_data; 
    end
    if(_T_user__T_10_en & _T_user__T_10_mask) begin
      _T_user[_T_user__T_10_addr] <= _T_user__T_10_data; 
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_3) begin
          if (io_deq_ready) begin
            _T_1 <= 1'h0;
          end else begin
            _T_1 <= _T_6;
          end
        end else begin
          _T_1 <= _T_6;
        end
      end
    end
  end
endmodule
module dual_Queue_67( 
  input        clock, 
  input        reset, 
  output       io_enq_ready, 
  input        io_enq_valid, 
  input  [2:0] io_enq_bits_opcode, 
  input  [2:0] io_enq_bits_size, 
  input  [6:0] io_enq_bits_source, 
  input        io_deq_ready, 
  output       io_deq_valid, 
  output [2:0] io_deq_bits_opcode, 
  output [2:0] io_deq_bits_size, 
  output [6:0] io_deq_bits_source 
);
  reg [2:0] _T_opcode [0:0]; 
  reg [31:0] _RAND_0;
  wire [2:0] _T_opcode__T_14_data; 
  wire  _T_opcode__T_14_addr; 
  wire [2:0] _T_opcode__T_10_data; 
  wire  _T_opcode__T_10_addr; 
  wire  _T_opcode__T_10_mask; 
  wire  _T_opcode__T_10_en; 
  reg [2:0] _T_size [0:0]; 
  reg [31:0] _RAND_1;
  wire [2:0] _T_size__T_14_data; 
  wire  _T_size__T_14_addr; 
  wire [2:0] _T_size__T_10_data; 
  wire  _T_size__T_10_addr; 
  wire  _T_size__T_10_mask; 
  wire  _T_size__T_10_en; 
  reg [6:0] _T_source [0:0]; 
  reg [31:0] _RAND_2;
  wire [6:0] _T_source__T_14_data; 
  wire  _T_source__T_14_addr; 
  wire [6:0] _T_source__T_10_data; 
  wire  _T_source__T_10_addr; 
  wire  _T_source__T_10_mask; 
  wire  _T_source__T_10_en; 
  reg  _T_1; 
  reg [31:0] _RAND_3;
  wire  _T_3; 
  wire  _T_6; 
  wire  _T_8; 
  wire  _T_11; 
  assign _T_opcode__T_14_addr = 1'h0;
  assign _T_opcode__T_14_data = _T_opcode[_T_opcode__T_14_addr]; 
  assign _T_opcode__T_10_data = io_enq_bits_opcode;
  assign _T_opcode__T_10_addr = 1'h0;
  assign _T_opcode__T_10_mask = 1'h1;
  assign _T_opcode__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_size__T_14_addr = 1'h0;
  assign _T_size__T_14_data = _T_size[_T_size__T_14_addr]; 
  assign _T_size__T_10_data = io_enq_bits_size;
  assign _T_size__T_10_addr = 1'h0;
  assign _T_size__T_10_mask = 1'h1;
  assign _T_size__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_source__T_14_addr = 1'h0;
  assign _T_source__T_14_data = _T_source[_T_source__T_14_addr]; 
  assign _T_source__T_10_data = io_enq_bits_source;
  assign _T_source__T_10_addr = 1'h0;
  assign _T_source__T_10_mask = 1'h1;
  assign _T_source__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _T_11 = _T_6 != _T_8; 
  assign io_enq_ready = _T_1 == 1'h0; 
  assign io_deq_valid = _T_3 == 1'h0; 
  assign io_deq_bits_opcode = _T_opcode__T_14_data; 
  assign io_deq_bits_size = _T_size__T_14_data; 
  assign io_deq_bits_source = _T_source__T_14_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_size[initvar] = _RAND_1[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_source[initvar] = _RAND_2[6:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T_opcode__T_10_en & _T_opcode__T_10_mask) begin
      _T_opcode[_T_opcode__T_10_addr] <= _T_opcode__T_10_data; 
    end
    if(_T_size__T_10_en & _T_size__T_10_mask) begin
      _T_size[_T_size__T_10_addr] <= _T_size__T_10_data; 
    end
    if(_T_source__T_10_en & _T_source__T_10_mask) begin
      _T_source[_T_source__T_10_addr] <= _T_source__T_10_data; 
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_11) begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module dual_Queue_68( 
  input        clock, 
  input        reset, 
  output       io_enq_ready, 
  input        io_enq_valid, 
  input  [2:0] io_enq_bits_opcode, 
  input  [2:0] io_enq_bits_param, 
  input  [2:0] io_enq_bits_size, 
  input  [6:0] io_enq_bits_source, 
  input        io_deq_ready, 
  output       io_deq_valid, 
  output [2:0] io_deq_bits_opcode, 
  output [2:0] io_deq_bits_param, 
  output [2:0] io_deq_bits_size, 
  output [6:0] io_deq_bits_source 
);
  reg [2:0] _T_opcode [0:0]; 
  reg [31:0] _RAND_0;
  wire [2:0] _T_opcode__T_14_data; 
  wire  _T_opcode__T_14_addr; 
  wire [2:0] _T_opcode__T_10_data; 
  wire  _T_opcode__T_10_addr; 
  wire  _T_opcode__T_10_mask; 
  wire  _T_opcode__T_10_en; 
  reg [2:0] _T_param [0:0]; 
  reg [31:0] _RAND_1;
  wire [2:0] _T_param__T_14_data; 
  wire  _T_param__T_14_addr; 
  wire [2:0] _T_param__T_10_data; 
  wire  _T_param__T_10_addr; 
  wire  _T_param__T_10_mask; 
  wire  _T_param__T_10_en; 
  reg [2:0] _T_size [0:0]; 
  reg [31:0] _RAND_2;
  wire [2:0] _T_size__T_14_data; 
  wire  _T_size__T_14_addr; 
  wire [2:0] _T_size__T_10_data; 
  wire  _T_size__T_10_addr; 
  wire  _T_size__T_10_mask; 
  wire  _T_size__T_10_en; 
  reg [6:0] _T_source [0:0]; 
  reg [31:0] _RAND_3;
  wire [6:0] _T_source__T_14_data; 
  wire  _T_source__T_14_addr; 
  wire [6:0] _T_source__T_10_data; 
  wire  _T_source__T_10_addr; 
  wire  _T_source__T_10_mask; 
  wire  _T_source__T_10_en; 
  reg  _T_1; 
  reg [31:0] _RAND_4;
  wire  _T_3; 
  wire  _T_6; 
  wire  _T_8; 
  wire  _T_11; 
  assign _T_opcode__T_14_addr = 1'h0;
  assign _T_opcode__T_14_data = _T_opcode[_T_opcode__T_14_addr]; 
  assign _T_opcode__T_10_data = io_enq_bits_opcode;
  assign _T_opcode__T_10_addr = 1'h0;
  assign _T_opcode__T_10_mask = 1'h1;
  assign _T_opcode__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_param__T_14_addr = 1'h0;
  assign _T_param__T_14_data = _T_param[_T_param__T_14_addr]; 
  assign _T_param__T_10_data = io_enq_bits_param;
  assign _T_param__T_10_addr = 1'h0;
  assign _T_param__T_10_mask = 1'h1;
  assign _T_param__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_size__T_14_addr = 1'h0;
  assign _T_size__T_14_data = _T_size[_T_size__T_14_addr]; 
  assign _T_size__T_10_data = io_enq_bits_size;
  assign _T_size__T_10_addr = 1'h0;
  assign _T_size__T_10_mask = 1'h1;
  assign _T_size__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_source__T_14_addr = 1'h0;
  assign _T_source__T_14_data = _T_source[_T_source__T_14_addr]; 
  assign _T_source__T_10_data = io_enq_bits_source;
  assign _T_source__T_10_addr = 1'h0;
  assign _T_source__T_10_mask = 1'h1;
  assign _T_source__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _T_11 = _T_6 != _T_8; 
  assign io_enq_ready = _T_1 == 1'h0; 
  assign io_deq_valid = _T_3 == 1'h0; 
  assign io_deq_bits_opcode = _T_opcode__T_14_data; 
  assign io_deq_bits_param = _T_param__T_14_data; 
  assign io_deq_bits_size = _T_size__T_14_data; 
  assign io_deq_bits_source = _T_source__T_14_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_param[initvar] = _RAND_1[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_size[initvar] = _RAND_2[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_source[initvar] = _RAND_3[6:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T_opcode__T_10_en & _T_opcode__T_10_mask) begin
      _T_opcode[_T_opcode__T_10_addr] <= _T_opcode__T_10_data; 
    end
    if(_T_param__T_10_en & _T_param__T_10_mask) begin
      _T_param[_T_param__T_10_addr] <= _T_param__T_10_data; 
    end
    if(_T_size__T_10_en & _T_size__T_10_mask) begin
      _T_size[_T_size__T_10_addr] <= _T_size__T_10_data; 
    end
    if(_T_source__T_10_en & _T_source__T_10_mask) begin
      _T_source[_T_source__T_10_addr] <= _T_source__T_10_data; 
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_11) begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module dual_Queue_8( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [2:0]  io_enq_bits_opcode, 
  input  [1:0]  io_enq_bits_param, 
  input  [3:0]  io_enq_bits_size, 
  input  [5:0]  io_enq_bits_source, 
  input         io_enq_bits_sink, 
  input         io_enq_bits_denied, 
  input  [31:0] io_enq_bits_data, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [2:0]  io_deq_bits_opcode, 
  output [1:0]  io_deq_bits_param, 
  output [3:0]  io_deq_bits_size, 
  output [5:0]  io_deq_bits_source, 
  output        io_deq_bits_sink, 
  output        io_deq_bits_denied, 
  output [31:0] io_deq_bits_data 
);
  reg [2:0] _T_opcode [0:0]; 
  reg [31:0] _RAND_0;
  wire [2:0] _T_opcode__T_14_data; 
  wire  _T_opcode__T_14_addr; 
  wire [2:0] _T_opcode__T_10_data; 
  wire  _T_opcode__T_10_addr; 
  wire  _T_opcode__T_10_mask; 
  wire  _T_opcode__T_10_en; 
  reg [1:0] _T_param [0:0]; 
  reg [31:0] _RAND_1;
  wire [1:0] _T_param__T_14_data; 
  wire  _T_param__T_14_addr; 
  wire [1:0] _T_param__T_10_data; 
  wire  _T_param__T_10_addr; 
  wire  _T_param__T_10_mask; 
  wire  _T_param__T_10_en; 
  reg [3:0] _T_size [0:0]; 
  reg [31:0] _RAND_2;
  wire [3:0] _T_size__T_14_data; 
  wire  _T_size__T_14_addr; 
  wire [3:0] _T_size__T_10_data; 
  wire  _T_size__T_10_addr; 
  wire  _T_size__T_10_mask; 
  wire  _T_size__T_10_en; 
  reg [5:0] _T_source [0:0]; 
  reg [31:0] _RAND_3;
  wire [5:0] _T_source__T_14_data; 
  wire  _T_source__T_14_addr; 
  wire [5:0] _T_source__T_10_data; 
  wire  _T_source__T_10_addr; 
  wire  _T_source__T_10_mask; 
  wire  _T_source__T_10_en; 
  reg  _T_sink [0:0]; 
  reg [31:0] _RAND_4;
  wire  _T_sink__T_14_data; 
  wire  _T_sink__T_14_addr; 
  wire  _T_sink__T_10_data; 
  wire  _T_sink__T_10_addr; 
  wire  _T_sink__T_10_mask; 
  wire  _T_sink__T_10_en; 
  reg  _T_denied [0:0]; 
  reg [31:0] _RAND_5;
  wire  _T_denied__T_14_data; 
  wire  _T_denied__T_14_addr; 
  wire  _T_denied__T_10_data; 
  wire  _T_denied__T_10_addr; 
  wire  _T_denied__T_10_mask; 
  wire  _T_denied__T_10_en; 
  reg [31:0] _T_data [0:0]; 
  reg [31:0] _RAND_6;
  wire [31:0] _T_data__T_14_data; 
  wire  _T_data__T_14_addr; 
  wire [31:0] _T_data__T_10_data; 
  wire  _T_data__T_10_addr; 
  wire  _T_data__T_10_mask; 
  wire  _T_data__T_10_en; 
  reg  _T_1; 
  reg [31:0] _RAND_7;
  wire  _T_3; 
  wire  _T_6; 
  wire  _T_8; 
  wire  _GEN_14; 
  wire  _GEN_24; 
  wire  _GEN_23; 
  wire  _T_11; 
  wire  _T_12; 
  assign _T_opcode__T_14_addr = 1'h0;
  assign _T_opcode__T_14_data = _T_opcode[_T_opcode__T_14_addr]; 
  assign _T_opcode__T_10_data = io_enq_bits_opcode;
  assign _T_opcode__T_10_addr = 1'h0;
  assign _T_opcode__T_10_mask = 1'h1;
  assign _T_opcode__T_10_en = _T_3 ? _GEN_14 : _T_6;
  assign _T_param__T_14_addr = 1'h0;
  assign _T_param__T_14_data = _T_param[_T_param__T_14_addr]; 
  assign _T_param__T_10_data = io_enq_bits_param;
  assign _T_param__T_10_addr = 1'h0;
  assign _T_param__T_10_mask = 1'h1;
  assign _T_param__T_10_en = _T_3 ? _GEN_14 : _T_6;
  assign _T_size__T_14_addr = 1'h0;
  assign _T_size__T_14_data = _T_size[_T_size__T_14_addr]; 
  assign _T_size__T_10_data = io_enq_bits_size;
  assign _T_size__T_10_addr = 1'h0;
  assign _T_size__T_10_mask = 1'h1;
  assign _T_size__T_10_en = _T_3 ? _GEN_14 : _T_6;
  assign _T_source__T_14_addr = 1'h0;
  assign _T_source__T_14_data = _T_source[_T_source__T_14_addr]; 
  assign _T_source__T_10_data = io_enq_bits_source;
  assign _T_source__T_10_addr = 1'h0;
  assign _T_source__T_10_mask = 1'h1;
  assign _T_source__T_10_en = _T_3 ? _GEN_14 : _T_6;
  assign _T_sink__T_14_addr = 1'h0;
  assign _T_sink__T_14_data = _T_sink[_T_sink__T_14_addr]; 
  assign _T_sink__T_10_data = io_enq_bits_sink;
  assign _T_sink__T_10_addr = 1'h0;
  assign _T_sink__T_10_mask = 1'h1;
  assign _T_sink__T_10_en = _T_3 ? _GEN_14 : _T_6;
  assign _T_denied__T_14_addr = 1'h0;
  assign _T_denied__T_14_data = _T_denied[_T_denied__T_14_addr]; 
  assign _T_denied__T_10_data = io_enq_bits_denied;
  assign _T_denied__T_10_addr = 1'h0;
  assign _T_denied__T_10_mask = 1'h1;
  assign _T_denied__T_10_en = _T_3 ? _GEN_14 : _T_6;
  assign _T_data__T_14_addr = 1'h0;
  assign _T_data__T_14_data = _T_data[_T_data__T_14_addr]; 
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = 1'h0;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = _T_3 ? _GEN_14 : _T_6;
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _GEN_14 = io_deq_ready ? 1'h0 : _T_6; 
  assign _GEN_24 = _T_3 ? _GEN_14 : _T_6; 
  assign _GEN_23 = _T_3 ? 1'h0 : _T_8; 
  assign _T_11 = _GEN_24 != _GEN_23; 
  assign _T_12 = _T_3 == 1'h0; 
  assign io_enq_ready = _T_1 == 1'h0; 
  assign io_deq_valid = io_enq_valid ? 1'h1 : _T_12; 
  assign io_deq_bits_opcode = _T_3 ? io_enq_bits_opcode : _T_opcode__T_14_data; 
  assign io_deq_bits_param = _T_3 ? io_enq_bits_param : _T_param__T_14_data; 
  assign io_deq_bits_size = _T_3 ? io_enq_bits_size : _T_size__T_14_data; 
  assign io_deq_bits_source = _T_3 ? io_enq_bits_source : _T_source__T_14_data; 
  assign io_deq_bits_sink = _T_3 ? io_enq_bits_sink : _T_sink__T_14_data; 
  assign io_deq_bits_denied = _T_3 ? io_enq_bits_denied : _T_denied__T_14_data; 
  assign io_deq_bits_data = _T_3 ? io_enq_bits_data : _T_data__T_14_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_param[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_size[initvar] = _RAND_2[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_source[initvar] = _RAND_3[5:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_sink[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_denied[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_data[initvar] = _RAND_6[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_1 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T_opcode__T_10_en & _T_opcode__T_10_mask) begin
      _T_opcode[_T_opcode__T_10_addr] <= _T_opcode__T_10_data; 
    end
    if(_T_param__T_10_en & _T_param__T_10_mask) begin
      _T_param[_T_param__T_10_addr] <= _T_param__T_10_data; 
    end
    if(_T_size__T_10_en & _T_size__T_10_mask) begin
      _T_size[_T_size__T_10_addr] <= _T_size__T_10_data; 
    end
    if(_T_source__T_10_en & _T_source__T_10_mask) begin
      _T_source[_T_source__T_10_addr] <= _T_source__T_10_data; 
    end
    if(_T_sink__T_10_en & _T_sink__T_10_mask) begin
      _T_sink[_T_sink__T_10_addr] <= _T_sink__T_10_data; 
    end
    if(_T_denied__T_10_en & _T_denied__T_10_mask) begin
      _T_denied[_T_denied__T_10_addr] <= _T_denied__T_10_data; 
    end
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; 
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_3) begin
          if (io_deq_ready) begin
            _T_1 <= 1'h0;
          end else begin
            _T_1 <= _T_6;
          end
        end else begin
          _T_1 <= _T_6;
        end
      end
    end
  end
endmodule
module dual_Queue_9( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [31:0] io_enq_bits, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [31:0] io_deq_bits 
);
  reg [31:0] _T [0:0]; 
  reg [31:0] _RAND_0;
  wire [31:0] _T__T_14_data; 
  wire  _T__T_14_addr; 
  wire [31:0] _T__T_10_data; 
  wire  _T__T_10_addr; 
  wire  _T__T_10_mask; 
  wire  _T__T_10_en; 
  reg  _T_1; 
  reg [31:0] _RAND_1;
  wire  _T_3; 
  wire  _T_6; 
  wire  _T_8; 
  wire  _T_11; 
  assign _T__T_14_addr = 1'h0;
  assign _T__T_14_data = _T[_T__T_14_addr]; 
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = 1'h0;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _T_11 = _T_6 != _T_8; 
  assign io_enq_ready = io_deq_ready ? 1'h1 : _T_3; 
  assign io_deq_valid = _T_3 == 1'h0; 
  assign io_deq_bits = _T__T_14_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; 
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_11) begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module dual_Queue( 
  input        clock, 
  input        reset, 
  output       io_enq_ready, 
  input        io_enq_valid, 
  input  [2:0] io_enq_bits_opcode, 
  input  [2:0] io_enq_bits_size, 
  input  [2:0] io_enq_bits_source, 
  input        io_deq_ready, 
  output       io_deq_valid, 
  output [2:0] io_deq_bits_opcode, 
  output [2:0] io_deq_bits_size, 
  output [2:0] io_deq_bits_source 
);
  reg [2:0] _T_opcode [0:0]; 
  reg [31:0] _RAND_0;
  wire [2:0] _T_opcode__T_14_data; 
  wire  _T_opcode__T_14_addr; 
  wire [2:0] _T_opcode__T_10_data; 
  wire  _T_opcode__T_10_addr; 
  wire  _T_opcode__T_10_mask; 
  wire  _T_opcode__T_10_en; 
  reg [2:0] _T_size [0:0]; 
  reg [31:0] _RAND_1;
  wire [2:0] _T_size__T_14_data; 
  wire  _T_size__T_14_addr; 
  wire [2:0] _T_size__T_10_data; 
  wire  _T_size__T_10_addr; 
  wire  _T_size__T_10_mask; 
  wire  _T_size__T_10_en; 
  reg [2:0] _T_source [0:0]; 
  reg [31:0] _RAND_2;
  wire [2:0] _T_source__T_14_data; 
  wire  _T_source__T_14_addr; 
  wire [2:0] _T_source__T_10_data; 
  wire  _T_source__T_10_addr; 
  wire  _T_source__T_10_mask; 
  wire  _T_source__T_10_en; 
  reg  _T_1; 
  reg [31:0] _RAND_3;
  wire  _T_3; 
  wire  _T_6; 
  wire  _T_8; 
  wire  _T_11; 
  assign _T_opcode__T_14_addr = 1'h0;
  assign _T_opcode__T_14_data = _T_opcode[_T_opcode__T_14_addr]; 
  assign _T_opcode__T_10_data = io_enq_bits_opcode;
  assign _T_opcode__T_10_addr = 1'h0;
  assign _T_opcode__T_10_mask = 1'h1;
  assign _T_opcode__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_size__T_14_addr = 1'h0;
  assign _T_size__T_14_data = _T_size[_T_size__T_14_addr]; 
  assign _T_size__T_10_data = io_enq_bits_size;
  assign _T_size__T_10_addr = 1'h0;
  assign _T_size__T_10_mask = 1'h1;
  assign _T_size__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_source__T_14_addr = 1'h0;
  assign _T_source__T_14_data = _T_source[_T_source__T_14_addr]; 
  assign _T_source__T_10_data = io_enq_bits_source;
  assign _T_source__T_10_addr = 1'h0;
  assign _T_source__T_10_mask = 1'h1;
  assign _T_source__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_3 = _T_1 == 1'h0; 
  assign _T_6 = io_enq_ready & io_enq_valid; 
  assign _T_8 = io_deq_ready & io_deq_valid; 
  assign _T_11 = _T_6 != _T_8; 
  assign io_enq_ready = _T_1 == 1'h0; 
  assign io_deq_valid = _T_3 == 1'h0; 
  assign io_deq_bits_opcode = _T_opcode__T_14_data; 
  assign io_deq_bits_size = _T_size__T_14_data; 
  assign io_deq_bits_source = _T_source__T_14_data; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_size[initvar] = _RAND_1[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_source[initvar] = _RAND_2[2:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if(_T_opcode__T_10_en & _T_opcode__T_10_mask) begin
      _T_opcode[_T_opcode__T_10_addr] <= _T_opcode__T_10_data; 
    end
    if(_T_size__T_10_en & _T_size__T_10_mask) begin
      _T_size[_T_size__T_10_addr] <= _T_size__T_10_data; 
    end
    if(_T_source__T_10_en & _T_source__T_10_mask) begin
      _T_source[_T_source__T_10_addr] <= _T_source__T_10_data; 
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      if (_T_11) begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module dual_ram_ext(
  input W0_clk,
  input [10:0] W0_addr,
  input W0_en,
  input [31:0] W0_data,
  input R0_clk,
  input [10:0] R0_addr,
  input R0_en,
  output [31:0] R0_data
);

  reg reg_R0_ren;
  reg [10:0] reg_R0_addr;
  reg [31:0] dual_ram [2047:0];
  `ifdef RANDOMIZE_MEM_INIT
    integer initvar;
    initial begin
      #`RANDOMIZE_DELAY begin end
      for (initvar = 0; initvar < 2048; initvar = initvar+1)
        dual_ram[initvar] = {1 {$random}};
      reg_R0_addr = {1 {$random}};
    end
  `endif
  integer i;
  always @(posedge R0_clk)
    reg_R0_ren <= R0_en;
  always @(posedge R0_clk)
    if (R0_en) reg_R0_addr <= R0_addr;
  always @(posedge W0_clk)
    if (W0_en) begin
      dual_ram[W0_addr][31:0] <= W0_data[31:0];
    end
  `ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] R0_random;
  `ifdef RANDOMIZE_MEM_INIT
    initial begin
      #`RANDOMIZE_DELAY begin end
      R0_random = {$random};
      reg_R0_ren = R0_random[0];
    end
  `endif
  always @(posedge R0_clk) R0_random <= {$random};
  assign R0_data = reg_R0_ren ? dual_ram[reg_R0_addr] : R0_random[31:0];
  `else
  assign R0_data = dual_ram[reg_R0_addr];
  `endif

endmodule

module dual_ram(
  input  [10:0] R0_addr,
  input         R0_en,
  input         R0_clk,
  output [31:0] R0_data,
  input  [10:0] W0_addr,
  input         W0_en,
  input         W0_clk,
  input  [31:0] W0_data
);
  wire [10:0] ram_ext_R0_addr;
  wire  ram_ext_R0_en;
  wire  ram_ext_R0_clk;
  wire [31:0] ram_ext_R0_data;
  wire [10:0] ram_ext_W0_addr;
  wire  ram_ext_W0_en;
  wire  ram_ext_W0_clk;
  wire [31:0] ram_ext_W0_data;
  dual_ram_ext ram_ext (
    .R0_addr(ram_ext_R0_addr),
    .R0_en(ram_ext_R0_en),
    .R0_clk(ram_ext_R0_clk),
    .R0_data(ram_ext_R0_data),
    .W0_addr(ram_ext_W0_addr),
    .W0_en(ram_ext_W0_en),
    .W0_clk(ram_ext_W0_clk),
    .W0_data(ram_ext_W0_data)
  );
  assign ram_ext_R0_clk = R0_clk;
  assign ram_ext_R0_en = R0_en;
  assign ram_ext_R0_addr = R0_addr;
  assign R0_data = $unsigned(ram_ext_R0_data);
  assign ram_ext_W0_clk = W0_clk;
  assign ram_ext_W0_en = W0_en;
  assign ram_ext_W0_addr = W0_addr;
  assign ram_ext_W0_data = $unsigned(W0_data);
endmodule
module dual_Repeater_1( 
  input         clock, 
  input         reset, 
  input         io_repeat, 
  output        io_full, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [3:0]  io_enq_bits_size, 
  input  [5:0]  io_enq_bits_source, 
  input  [31:0] io_enq_bits_address, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [3:0]  io_deq_bits_size, 
  output [5:0]  io_deq_bits_source, 
  output [31:0] io_deq_bits_address 
);
  reg  full; 
  reg [31:0] _RAND_0;
  reg [3:0] saved_size; 
  reg [31:0] _RAND_1;
  reg [5:0] saved_source; 
  reg [31:0] _RAND_2;
  reg [31:0] saved_address; 
  reg [31:0] _RAND_3;
  wire  _T_1; 
  wire  _T_4; 
  wire  _T_5; 
  wire  _T_6; 
  wire  _T_7; 
  wire  _T_8; 
  assign _T_1 = full == 1'h0; 
  assign _T_4 = io_enq_ready & io_enq_valid; 
  assign _T_5 = _T_4 & io_repeat; 
  assign _T_6 = io_deq_ready & io_deq_valid; 
  assign _T_7 = io_repeat == 1'h0; 
  assign _T_8 = _T_6 & _T_7; 
  assign io_full = full; 
  assign io_enq_ready = io_deq_ready & _T_1; 
  assign io_deq_valid = io_enq_valid | full; 
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; 
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; 
  assign io_deq_bits_address = full ? saved_address : io_enq_bits_address; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  saved_size = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  saved_source = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  saved_address = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      full <= 1'h0;
    end else begin
      if (_T_8) begin
        full <= 1'h0;
      end else begin
        if (_T_5) begin
          full <= 1'h1;
        end
      end
    end
    if (_T_5) begin
      saved_size <= io_enq_bits_size;
    end
    if (_T_5) begin
      saved_source <= io_enq_bits_source;
    end
    if (_T_5) begin
      saved_address <= io_enq_bits_address;
    end
  end
endmodule
module dual_Repeater_2( 
  input         clock, 
  input         reset, 
  input         io_repeat, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [2:0]  io_enq_bits_opcode, 
  input  [1:0]  io_enq_bits_param, 
  input  [3:0]  io_enq_bits_size, 
  input  [5:0]  io_enq_bits_source, 
  input         io_enq_bits_sink, 
  input         io_enq_bits_denied, 
  input  [63:0] io_enq_bits_data, 
  input         io_enq_bits_corrupt, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [2:0]  io_deq_bits_opcode, 
  output [1:0]  io_deq_bits_param, 
  output [3:0]  io_deq_bits_size, 
  output [5:0]  io_deq_bits_source, 
  output        io_deq_bits_sink, 
  output        io_deq_bits_denied, 
  output [63:0] io_deq_bits_data, 
  output        io_deq_bits_corrupt 
);
  reg  full; 
  reg [31:0] _RAND_0;
  reg [2:0] saved_opcode; 
  reg [31:0] _RAND_1;
  reg [1:0] saved_param; 
  reg [31:0] _RAND_2;
  reg [3:0] saved_size; 
  reg [31:0] _RAND_3;
  reg [5:0] saved_source; 
  reg [31:0] _RAND_4;
  reg  saved_sink; 
  reg [31:0] _RAND_5;
  reg  saved_denied; 
  reg [31:0] _RAND_6;
  reg [63:0] saved_data; 
  reg [63:0] _RAND_7;
  reg  saved_corrupt; 
  reg [31:0] _RAND_8;
  wire  _T_1; 
  wire  _T_4; 
  wire  _T_5; 
  wire  _T_6; 
  wire  _T_7; 
  wire  _T_8; 
  assign _T_1 = full == 1'h0; 
  assign _T_4 = io_enq_ready & io_enq_valid; 
  assign _T_5 = _T_4 & io_repeat; 
  assign _T_6 = io_deq_ready & io_deq_valid; 
  assign _T_7 = io_repeat == 1'h0; 
  assign _T_8 = _T_6 & _T_7; 
  assign io_enq_ready = io_deq_ready & _T_1; 
  assign io_deq_valid = io_enq_valid | full; 
  assign io_deq_bits_opcode = full ? saved_opcode : io_enq_bits_opcode; 
  assign io_deq_bits_param = full ? saved_param : io_enq_bits_param; 
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; 
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; 
  assign io_deq_bits_sink = full ? saved_sink : io_enq_bits_sink; 
  assign io_deq_bits_denied = full ? saved_denied : io_enq_bits_denied; 
  assign io_deq_bits_data = full ? saved_data : io_enq_bits_data; 
  assign io_deq_bits_corrupt = full ? saved_corrupt : io_enq_bits_corrupt; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  saved_opcode = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  saved_param = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  saved_size = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  saved_source = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  saved_sink = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  saved_denied = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{`RANDOM}};
  saved_data = _RAND_7[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  saved_corrupt = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      full <= 1'h0;
    end else begin
      if (_T_8) begin
        full <= 1'h0;
      end else begin
        if (_T_5) begin
          full <= 1'h1;
        end
      end
    end
    if (_T_5) begin
      saved_opcode <= io_enq_bits_opcode;
    end
    if (_T_5) begin
      saved_param <= io_enq_bits_param;
    end
    if (_T_5) begin
      saved_size <= io_enq_bits_size;
    end
    if (_T_5) begin
      saved_source <= io_enq_bits_source;
    end
    if (_T_5) begin
      saved_sink <= io_enq_bits_sink;
    end
    if (_T_5) begin
      saved_denied <= io_enq_bits_denied;
    end
    if (_T_5) begin
      saved_data <= io_enq_bits_data;
    end
    if (_T_5) begin
      saved_corrupt <= io_enq_bits_corrupt;
    end
  end
endmodule
module dual_Repeater_4( 
  input         clock, 
  input         reset, 
  input         io_repeat, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [2:0]  io_enq_bits_opcode, 
  input  [2:0]  io_enq_bits_param, 
  input  [2:0]  io_enq_bits_size, 
  input  [6:0]  io_enq_bits_source, 
  input  [28:0] io_enq_bits_address, 
  input  [7:0]  io_enq_bits_mask, 
  input         io_enq_bits_corrupt, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [2:0]  io_deq_bits_opcode, 
  output [2:0]  io_deq_bits_param, 
  output [2:0]  io_deq_bits_size, 
  output [6:0]  io_deq_bits_source, 
  output [28:0] io_deq_bits_address, 
  output [7:0]  io_deq_bits_mask, 
  output        io_deq_bits_corrupt 
);
  reg  full; 
  reg [31:0] _RAND_0;
  reg [2:0] saved_opcode; 
  reg [31:0] _RAND_1;
  reg [2:0] saved_param; 
  reg [31:0] _RAND_2;
  reg [2:0] saved_size; 
  reg [31:0] _RAND_3;
  reg [6:0] saved_source; 
  reg [31:0] _RAND_4;
  reg [28:0] saved_address; 
  reg [31:0] _RAND_5;
  reg [7:0] saved_mask; 
  reg [31:0] _RAND_6;
  reg  saved_corrupt; 
  reg [31:0] _RAND_7;
  wire  _T_1; 
  wire  _T_4; 
  wire  _T_5; 
  wire  _T_6; 
  wire  _T_7; 
  wire  _T_8; 
  assign _T_1 = full == 1'h0; 
  assign _T_4 = io_enq_ready & io_enq_valid; 
  assign _T_5 = _T_4 & io_repeat; 
  assign _T_6 = io_deq_ready & io_deq_valid; 
  assign _T_7 = io_repeat == 1'h0; 
  assign _T_8 = _T_6 & _T_7; 
  assign io_enq_ready = io_deq_ready & _T_1; 
  assign io_deq_valid = io_enq_valid | full; 
  assign io_deq_bits_opcode = full ? saved_opcode : io_enq_bits_opcode; 
  assign io_deq_bits_param = full ? saved_param : io_enq_bits_param; 
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; 
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; 
  assign io_deq_bits_address = full ? saved_address : io_enq_bits_address; 
  assign io_deq_bits_mask = full ? saved_mask : io_enq_bits_mask; 
  assign io_deq_bits_corrupt = full ? saved_corrupt : io_enq_bits_corrupt; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  saved_opcode = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  saved_param = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  saved_size = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  saved_source = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  saved_address = _RAND_5[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  saved_mask = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  saved_corrupt = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      full <= 1'h0;
    end else begin
      if (_T_8) begin
        full <= 1'h0;
      end else begin
        if (_T_5) begin
          full <= 1'h1;
        end
      end
    end
    if (_T_5) begin
      saved_opcode <= io_enq_bits_opcode;
    end
    if (_T_5) begin
      saved_param <= io_enq_bits_param;
    end
    if (_T_5) begin
      saved_size <= io_enq_bits_size;
    end
    if (_T_5) begin
      saved_source <= io_enq_bits_source;
    end
    if (_T_5) begin
      saved_address <= io_enq_bits_address;
    end
    if (_T_5) begin
      saved_mask <= io_enq_bits_mask;
    end
    if (_T_5) begin
      saved_corrupt <= io_enq_bits_corrupt;
    end
  end
endmodule
module dual_Repeater_5( 
  input         clock, 
  input         reset, 
  input         io_repeat, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [2:0]  io_enq_bits_opcode, 
  input  [2:0]  io_enq_bits_param, 
  input  [2:0]  io_enq_bits_size, 
  input  [6:0]  io_enq_bits_source, 
  input  [28:0] io_enq_bits_address, 
  input         io_enq_bits_corrupt, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [2:0]  io_deq_bits_opcode, 
  output [2:0]  io_deq_bits_param, 
  output [2:0]  io_deq_bits_size, 
  output [6:0]  io_deq_bits_source, 
  output [28:0] io_deq_bits_address, 
  output        io_deq_bits_corrupt 
);
  reg  full; 
  reg [31:0] _RAND_0;
  reg [2:0] saved_opcode; 
  reg [31:0] _RAND_1;
  reg [2:0] saved_param; 
  reg [31:0] _RAND_2;
  reg [2:0] saved_size; 
  reg [31:0] _RAND_3;
  reg [6:0] saved_source; 
  reg [31:0] _RAND_4;
  reg [28:0] saved_address; 
  reg [31:0] _RAND_5;
  reg  saved_corrupt; 
  reg [31:0] _RAND_6;
  wire  _T_1; 
  wire  _T_4; 
  wire  _T_5; 
  wire  _T_6; 
  wire  _T_7; 
  wire  _T_8; 
  assign _T_1 = full == 1'h0; 
  assign _T_4 = io_enq_ready & io_enq_valid; 
  assign _T_5 = _T_4 & io_repeat; 
  assign _T_6 = io_deq_ready & io_deq_valid; 
  assign _T_7 = io_repeat == 1'h0; 
  assign _T_8 = _T_6 & _T_7; 
  assign io_enq_ready = io_deq_ready & _T_1; 
  assign io_deq_valid = io_enq_valid | full; 
  assign io_deq_bits_opcode = full ? saved_opcode : io_enq_bits_opcode; 
  assign io_deq_bits_param = full ? saved_param : io_enq_bits_param; 
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; 
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; 
  assign io_deq_bits_address = full ? saved_address : io_enq_bits_address; 
  assign io_deq_bits_corrupt = full ? saved_corrupt : io_enq_bits_corrupt; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  saved_opcode = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  saved_param = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  saved_size = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  saved_source = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  saved_address = _RAND_5[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  saved_corrupt = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      full <= 1'h0;
    end else begin
      if (_T_8) begin
        full <= 1'h0;
      end else begin
        if (_T_5) begin
          full <= 1'h1;
        end
      end
    end
    if (_T_5) begin
      saved_opcode <= io_enq_bits_opcode;
    end
    if (_T_5) begin
      saved_param <= io_enq_bits_param;
    end
    if (_T_5) begin
      saved_size <= io_enq_bits_size;
    end
    if (_T_5) begin
      saved_source <= io_enq_bits_source;
    end
    if (_T_5) begin
      saved_address <= io_enq_bits_address;
    end
    if (_T_5) begin
      saved_corrupt <= io_enq_bits_corrupt;
    end
  end
endmodule
module dual_Repeater_top( 
  input         clock, 
  input         reset, 
  input         io_repeat, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [2:0]  io_enq_bits_opcode, 
  input  [2:0]  io_enq_bits_param, 
  input  [2:0]  io_enq_bits_size, 
  input  [2:0]  io_enq_bits_source, 
  input  [31:0] io_enq_bits_address, 
  input  [7:0]  io_enq_bits_mask, 
  input  [63:0] io_enq_bits_data, 
  input         io_enq_bits_corrupt, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [2:0]  io_deq_bits_opcode, 
  output [2:0]  io_deq_bits_param, 
  output [2:0]  io_deq_bits_size, 
  output [2:0]  io_deq_bits_source, 
  output [31:0] io_deq_bits_address, 
  output [7:0]  io_deq_bits_mask, 
  output [63:0] io_deq_bits_data, 
  output        io_deq_bits_corrupt 
);
  reg  full; 
  reg [31:0] _RAND_0;
  reg [2:0] saved_opcode; 
  reg [31:0] _RAND_1;
  reg [2:0] saved_param; 
  reg [31:0] _RAND_2;
  reg [2:0] saved_size; 
  reg [31:0] _RAND_3;
  reg [2:0] saved_source; 
  reg [31:0] _RAND_4;
  reg [31:0] saved_address; 
  reg [31:0] _RAND_5;
  reg [7:0] saved_mask; 
  reg [31:0] _RAND_6;
  reg [63:0] saved_data; 
  reg [63:0] _RAND_7;
  reg  saved_corrupt; 
  reg [31:0] _RAND_8;
  wire  _T_1; 
  wire  _T_4; 
  wire  _T_5; 
  wire  _T_6; 
  wire  _T_7; 
  wire  _T_8; 
  assign _T_1 = full == 1'h0; 
  assign _T_4 = io_enq_ready & io_enq_valid; 
  assign _T_5 = _T_4 & io_repeat; 
  assign _T_6 = io_deq_ready & io_deq_valid; 
  assign _T_7 = io_repeat == 1'h0; 
  assign _T_8 = _T_6 & _T_7; 
  assign io_enq_ready = io_deq_ready & _T_1; 
  assign io_deq_valid = io_enq_valid | full; 
  assign io_deq_bits_opcode = full ? saved_opcode : io_enq_bits_opcode; 
  assign io_deq_bits_param = full ? saved_param : io_enq_bits_param; 
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; 
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; 
  assign io_deq_bits_address = full ? saved_address : io_enq_bits_address; 
  assign io_deq_bits_mask = full ? saved_mask : io_enq_bits_mask; 
  assign io_deq_bits_data = full ? saved_data : io_enq_bits_data; 
  assign io_deq_bits_corrupt = full ? saved_corrupt : io_enq_bits_corrupt; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  saved_opcode = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  saved_param = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  saved_size = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  saved_source = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  saved_address = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  saved_mask = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{`RANDOM}};
  saved_data = _RAND_7[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  saved_corrupt = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      full <= 1'h0;
    end else begin
      if (_T_8) begin
        full <= 1'h0;
      end else begin
        if (_T_5) begin
          full <= 1'h1;
        end
      end
    end
    if (_T_5) begin
      saved_opcode <= io_enq_bits_opcode;
    end
    if (_T_5) begin
      saved_param <= io_enq_bits_param;
    end
    if (_T_5) begin
      saved_size <= io_enq_bits_size;
    end
    if (_T_5) begin
      saved_source <= io_enq_bits_source;
    end
    if (_T_5) begin
      saved_address <= io_enq_bits_address;
    end
    if (_T_5) begin
      saved_mask <= io_enq_bits_mask;
    end
    if (_T_5) begin
      saved_data <= io_enq_bits_data;
    end
    if (_T_5) begin
      saved_corrupt <= io_enq_bits_corrupt;
    end
  end
endmodule
module dual_ResetCatchAndSync_d3( 
  input   clock, 
  input   reset, 
  output  io_sync_reset 
);
  wire  AsyncResetSynchronizerShiftReg_w1_d3_i0_clock; 
  wire  AsyncResetSynchronizerShiftReg_w1_d3_i0_reset; 
  wire  AsyncResetSynchronizerShiftReg_w1_d3_i0_io_d; 
  wire  AsyncResetSynchronizerShiftReg_w1_d3_i0_io_q; 
  wire  _T; 
  dual_AsyncResetSynchronizerShiftReg_w1_d3_i0 AsyncResetSynchronizerShiftReg_w1_d3_i0 ( 
    .clock(AsyncResetSynchronizerShiftReg_w1_d3_i0_clock),
    .reset(AsyncResetSynchronizerShiftReg_w1_d3_i0_reset),
    .io_d(AsyncResetSynchronizerShiftReg_w1_d3_i0_io_d),
    .io_q(AsyncResetSynchronizerShiftReg_w1_d3_i0_io_q)
  );
  assign _T = AsyncResetSynchronizerShiftReg_w1_d3_i0_io_q; 
  assign io_sync_reset = ~ _T; 
  assign AsyncResetSynchronizerShiftReg_w1_d3_i0_clock = clock; 
  assign AsyncResetSynchronizerShiftReg_w1_d3_i0_reset = reset; 
  assign AsyncResetSynchronizerShiftReg_w1_d3_i0_io_d = 1'h1; 
endmodule
module dual_RX( 
  input         clock, 
  input         reset, 
  input         io_b2c_send, 
  input  [31:0] io_b2c_data, 
  output [31:0] io_a_mem_0, 
  output [31:0] io_a_mem_1, 
  output [31:0] io_a_mem_2, 
  output [31:0] io_a_mem_3, 
  output [31:0] io_a_mem_4, 
  output [31:0] io_a_mem_5, 
  output [31:0] io_a_mem_6, 
  output [31:0] io_a_mem_7, 
  input  [3:0]  io_a_ridx, 
  output [3:0]  io_a_widx, 
  input         io_a_safe_ridx_valid, 
  output        io_a_safe_widx_valid, 
  output        io_a_safe_source_reset_n, 
  input         io_a_safe_sink_reset_n, 
  output [31:0] io_bmem_0, 
  output [31:0] io_bmem_1, 
  output [31:0] io_bmem_2, 
  output [31:0] io_bmem_3, 
  output [31:0] io_bmem_4, 
  output [31:0] io_bmem_5, 
  output [31:0] io_bmem_6, 
  output [31:0] io_bmem_7, 
  input  [3:0]  io_bridx, 
  output [3:0]  io_bwidx, 
  input         io_bsafe_ridx_valid, 
  output        io_bsafe_widx_valid, 
  output        io_bsafe_source_reset_n, 
  input         io_bsafe_sink_reset_n, 
  output [31:0] io_c_mem_0, 
  output [31:0] io_c_mem_1, 
  output [31:0] io_c_mem_2, 
  output [31:0] io_c_mem_3, 
  output [31:0] io_c_mem_4, 
  output [31:0] io_c_mem_5, 
  output [31:0] io_c_mem_6, 
  output [31:0] io_c_mem_7, 
  input  [3:0]  io_c_ridx, 
  output [3:0]  io_c_widx, 
  input         io_c_safe_ridx_valid, 
  output        io_c_safe_widx_valid, 
  output        io_c_safe_source_reset_n, 
  input         io_c_safe_sink_reset_n, 
  output [31:0] io_d_mem_0, 
  output [31:0] io_d_mem_1, 
  output [31:0] io_d_mem_2, 
  output [31:0] io_d_mem_3, 
  output [31:0] io_d_mem_4, 
  output [31:0] io_d_mem_5, 
  output [31:0] io_d_mem_6, 
  output [31:0] io_d_mem_7, 
  input  [3:0]  io_d_ridx, 
  output [3:0]  io_d_widx, 
  input         io_d_safe_ridx_valid, 
  output        io_d_safe_widx_valid, 
  output        io_d_safe_source_reset_n, 
  input         io_d_safe_sink_reset_n, 
  output [31:0] io_e_mem_0, 
  output [31:0] io_e_mem_1, 
  output [31:0] io_e_mem_2, 
  output [31:0] io_e_mem_3, 
  output [31:0] io_e_mem_4, 
  output [31:0] io_e_mem_5, 
  output [31:0] io_e_mem_6, 
  output [31:0] io_e_mem_7, 
  input  [3:0]  io_e_ridx, 
  output [3:0]  io_e_widx, 
  input         io_e_safe_ridx_valid, 
  output        io_e_safe_widx_valid, 
  output        io_e_safe_source_reset_n, 
  input         io_e_safe_sink_reset_n, 
  output [19:0] io_rxc_mem_0_a, 
  output [19:0] io_rxc_mem_0_b, 
  output [19:0] io_rxc_mem_0_c, 
  output [19:0] io_rxc_mem_0_d, 
  output [19:0] io_rxc_mem_0_e, 
  input         io_rxc_ridx, 
  output        io_rxc_widx, 
  input         io_rxc_safe_ridx_valid, 
  output        io_rxc_safe_widx_valid, 
  output        io_rxc_safe_source_reset_n, 
  input         io_rxc_safe_sink_reset_n, 
  output [19:0] io_txc_mem_0_a, 
  output [19:0] io_txc_mem_0_b, 
  output [19:0] io_txc_mem_0_c, 
  output [19:0] io_txc_mem_0_d, 
  output [19:0] io_txc_mem_0_e, 
  input         io_txc_ridx, 
  output        io_txc_widx, 
  input         io_txc_safe_ridx_valid, 
  output        io_txc_safe_widx_valid, 
  output        io_txc_safe_source_reset_n, 
  input         io_txc_safe_sink_reset_n 
);
  wire  hqa_clock; 
  wire  hqa_reset; 
  wire  hqa_io_enq_ready; 
  wire  hqa_io_enq_valid; 
  wire [31:0] hqa_io_enq_bits; 
  wire  hqa_io_deq_ready; 
  wire  hqa_io_deq_valid; 
  wire [31:0] hqa_io_deq_bits; 
  wire  hqb_clock; 
  wire  hqb_reset; 
  wire  hqb_io_enq_ready; 
  wire  hqb_io_enq_valid; 
  wire [31:0] hqb_io_enq_bits; 
  wire  hqb_io_deq_ready; 
  wire  hqb_io_deq_valid; 
  wire [31:0] hqb_io_deq_bits; 
  wire  hqc_clock; 
  wire  hqc_reset; 
  wire  hqc_io_enq_ready; 
  wire  hqc_io_enq_valid; 
  wire [31:0] hqc_io_enq_bits; 
  wire  hqc_io_deq_ready; 
  wire  hqc_io_deq_valid; 
  wire [31:0] hqc_io_deq_bits; 
  wire  hqd_clock; 
  wire  hqd_reset; 
  wire  hqd_io_enq_ready; 
  wire  hqd_io_enq_valid; 
  wire [31:0] hqd_io_enq_bits; 
  wire  hqd_io_deq_ready; 
  wire  hqd_io_deq_valid; 
  wire [31:0] hqd_io_deq_bits; 
  wire  hqe_clock; 
  wire  hqe_reset; 
  wire  hqe_io_enq_ready; 
  wire  hqe_io_enq_valid; 
  wire [31:0] hqe_io_enq_bits; 
  wire  hqe_io_deq_ready; 
  wire  hqe_io_deq_valid; 
  wire [31:0] hqe_io_deq_bits; 
  wire  AsyncQueueSource_clock; 
  wire  AsyncQueueSource_reset; 
  wire  AsyncQueueSource_io_enq_ready; 
  wire  AsyncQueueSource_io_enq_valid; 
  wire [31:0] AsyncQueueSource_io_enq_bits; 
  wire [31:0] AsyncQueueSource_io_async_mem_0; 
  wire [31:0] AsyncQueueSource_io_async_mem_1; 
  wire [31:0] AsyncQueueSource_io_async_mem_2; 
  wire [31:0] AsyncQueueSource_io_async_mem_3; 
  wire [31:0] AsyncQueueSource_io_async_mem_4; 
  wire [31:0] AsyncQueueSource_io_async_mem_5; 
  wire [31:0] AsyncQueueSource_io_async_mem_6; 
  wire [31:0] AsyncQueueSource_io_async_mem_7; 
  wire [3:0] AsyncQueueSource_io_async_ridx; 
  wire [3:0] AsyncQueueSource_io_async_widx; 
  wire  AsyncQueueSource_io_async_safe_ridx_valid; 
  wire  AsyncQueueSource_io_async_safe_widx_valid; 
  wire  AsyncQueueSource_io_async_safe_source_reset_n; 
  wire  AsyncQueueSource_io_async_safe_sink_reset_n; 
  wire  AsyncQueueSource_1_clock; 
  wire  AsyncQueueSource_1_reset; 
  wire  AsyncQueueSource_1_io_enq_ready; 
  wire  AsyncQueueSource_1_io_enq_valid; 
  wire [31:0] AsyncQueueSource_1_io_enq_bits; 
  wire [31:0] AsyncQueueSource_1_io_async_mem_0; 
  wire [31:0] AsyncQueueSource_1_io_async_mem_1; 
  wire [31:0] AsyncQueueSource_1_io_async_mem_2; 
  wire [31:0] AsyncQueueSource_1_io_async_mem_3; 
  wire [31:0] AsyncQueueSource_1_io_async_mem_4; 
  wire [31:0] AsyncQueueSource_1_io_async_mem_5; 
  wire [31:0] AsyncQueueSource_1_io_async_mem_6; 
  wire [31:0] AsyncQueueSource_1_io_async_mem_7; 
  wire [3:0] AsyncQueueSource_1_io_async_ridx; 
  wire [3:0] AsyncQueueSource_1_io_async_widx; 
  wire  AsyncQueueSource_1_io_async_safe_ridx_valid; 
  wire  AsyncQueueSource_1_io_async_safe_widx_valid; 
  wire  AsyncQueueSource_1_io_async_safe_source_reset_n; 
  wire  AsyncQueueSource_1_io_async_safe_sink_reset_n; 
  wire  AsyncQueueSource_2_clock; 
  wire  AsyncQueueSource_2_reset; 
  wire  AsyncQueueSource_2_io_enq_ready; 
  wire  AsyncQueueSource_2_io_enq_valid; 
  wire [31:0] AsyncQueueSource_2_io_enq_bits; 
  wire [31:0] AsyncQueueSource_2_io_async_mem_0; 
  wire [31:0] AsyncQueueSource_2_io_async_mem_1; 
  wire [31:0] AsyncQueueSource_2_io_async_mem_2; 
  wire [31:0] AsyncQueueSource_2_io_async_mem_3; 
  wire [31:0] AsyncQueueSource_2_io_async_mem_4; 
  wire [31:0] AsyncQueueSource_2_io_async_mem_5; 
  wire [31:0] AsyncQueueSource_2_io_async_mem_6; 
  wire [31:0] AsyncQueueSource_2_io_async_mem_7; 
  wire [3:0] AsyncQueueSource_2_io_async_ridx; 
  wire [3:0] AsyncQueueSource_2_io_async_widx; 
  wire  AsyncQueueSource_2_io_async_safe_ridx_valid; 
  wire  AsyncQueueSource_2_io_async_safe_widx_valid; 
  wire  AsyncQueueSource_2_io_async_safe_source_reset_n; 
  wire  AsyncQueueSource_2_io_async_safe_sink_reset_n; 
  wire  AsyncQueueSource_3_clock; 
  wire  AsyncQueueSource_3_reset; 
  wire  AsyncQueueSource_3_io_enq_ready; 
  wire  AsyncQueueSource_3_io_enq_valid; 
  wire [31:0] AsyncQueueSource_3_io_enq_bits; 
  wire [31:0] AsyncQueueSource_3_io_async_mem_0; 
  wire [31:0] AsyncQueueSource_3_io_async_mem_1; 
  wire [31:0] AsyncQueueSource_3_io_async_mem_2; 
  wire [31:0] AsyncQueueSource_3_io_async_mem_3; 
  wire [31:0] AsyncQueueSource_3_io_async_mem_4; 
  wire [31:0] AsyncQueueSource_3_io_async_mem_5; 
  wire [31:0] AsyncQueueSource_3_io_async_mem_6; 
  wire [31:0] AsyncQueueSource_3_io_async_mem_7; 
  wire [3:0] AsyncQueueSource_3_io_async_ridx; 
  wire [3:0] AsyncQueueSource_3_io_async_widx; 
  wire  AsyncQueueSource_3_io_async_safe_ridx_valid; 
  wire  AsyncQueueSource_3_io_async_safe_widx_valid; 
  wire  AsyncQueueSource_3_io_async_safe_source_reset_n; 
  wire  AsyncQueueSource_3_io_async_safe_sink_reset_n; 
  wire  AsyncQueueSource_4_clock; 
  wire  AsyncQueueSource_4_reset; 
  wire  AsyncQueueSource_4_io_enq_ready; 
  wire  AsyncQueueSource_4_io_enq_valid; 
  wire [31:0] AsyncQueueSource_4_io_enq_bits; 
  wire [31:0] AsyncQueueSource_4_io_async_mem_0; 
  wire [31:0] AsyncQueueSource_4_io_async_mem_1; 
  wire [31:0] AsyncQueueSource_4_io_async_mem_2; 
  wire [31:0] AsyncQueueSource_4_io_async_mem_3; 
  wire [31:0] AsyncQueueSource_4_io_async_mem_4; 
  wire [31:0] AsyncQueueSource_4_io_async_mem_5; 
  wire [31:0] AsyncQueueSource_4_io_async_mem_6; 
  wire [31:0] AsyncQueueSource_4_io_async_mem_7; 
  wire [3:0] AsyncQueueSource_4_io_async_ridx; 
  wire [3:0] AsyncQueueSource_4_io_async_widx; 
  wire  AsyncQueueSource_4_io_async_safe_ridx_valid; 
  wire  AsyncQueueSource_4_io_async_safe_widx_valid; 
  wire  AsyncQueueSource_4_io_async_safe_source_reset_n; 
  wire  AsyncQueueSource_4_io_async_safe_sink_reset_n; 
  wire  AsyncQueueSource_5_clock; 
  wire  AsyncQueueSource_5_reset; 
  wire  AsyncQueueSource_5_io_enq_ready; 
  wire  AsyncQueueSource_5_io_enq_valid; 
  wire [19:0] AsyncQueueSource_5_io_enq_bits_a; 
  wire [19:0] AsyncQueueSource_5_io_enq_bits_b; 
  wire [19:0] AsyncQueueSource_5_io_enq_bits_c; 
  wire [19:0] AsyncQueueSource_5_io_enq_bits_d; 
  wire [19:0] AsyncQueueSource_5_io_enq_bits_e; 
  wire [19:0] AsyncQueueSource_5_io_async_mem_0_a; 
  wire [19:0] AsyncQueueSource_5_io_async_mem_0_b; 
  wire [19:0] AsyncQueueSource_5_io_async_mem_0_c; 
  wire [19:0] AsyncQueueSource_5_io_async_mem_0_d; 
  wire [19:0] AsyncQueueSource_5_io_async_mem_0_e; 
  wire  AsyncQueueSource_5_io_async_ridx; 
  wire  AsyncQueueSource_5_io_async_widx; 
  wire  AsyncQueueSource_5_io_async_safe_ridx_valid; 
  wire  AsyncQueueSource_5_io_async_safe_widx_valid; 
  wire  AsyncQueueSource_5_io_async_safe_source_reset_n; 
  wire  AsyncQueueSource_5_io_async_safe_sink_reset_n; 
  wire  AsyncQueueSource_6_clock; 
  wire  AsyncQueueSource_6_reset; 
  wire  AsyncQueueSource_6_io_enq_ready; 
  wire  AsyncQueueSource_6_io_enq_valid; 
  wire [19:0] AsyncQueueSource_6_io_enq_bits_a; 
  wire [19:0] AsyncQueueSource_6_io_enq_bits_b; 
  wire [19:0] AsyncQueueSource_6_io_enq_bits_c; 
  wire [19:0] AsyncQueueSource_6_io_enq_bits_d; 
  wire [19:0] AsyncQueueSource_6_io_enq_bits_e; 
  wire [19:0] AsyncQueueSource_6_io_async_mem_0_a; 
  wire [19:0] AsyncQueueSource_6_io_async_mem_0_b; 
  wire [19:0] AsyncQueueSource_6_io_async_mem_0_c; 
  wire [19:0] AsyncQueueSource_6_io_async_mem_0_d; 
  wire [19:0] AsyncQueueSource_6_io_async_mem_0_e; 
  wire  AsyncQueueSource_6_io_async_ridx; 
  wire  AsyncQueueSource_6_io_async_widx; 
  wire  AsyncQueueSource_6_io_async_safe_ridx_valid; 
  wire  AsyncQueueSource_6_io_async_safe_widx_valid; 
  wire  AsyncQueueSource_6_io_async_safe_source_reset_n; 
  wire  AsyncQueueSource_6_io_async_safe_sink_reset_n; 
  reg [31:0] _T; 
  reg [31:0] _RAND_0;
  reg [31:0] b2c_data; 
  reg [31:0] _RAND_1;
  reg  _T_1; 
  reg [31:0] _RAND_2;
  reg  b2c_send; 
  reg [31:0] _RAND_3;
  reg [10:0] _T_2; 
  reg [31:0] _RAND_4;
  wire [2:0] _T_3; 
  wire [2:0] _T_4; 
  wire [3:0] _T_6; 
  wire [15:0] _T_11; 
  wire [12:0] _T_12; 
  wire [9:0] _T_13; 
  wire  _T_14; 
  wire [10:0] _T_15; 
  wire [6:0] _T_20; 
  wire  _T_21; 
  wire [7:0] _T_22; 
  wire  _T_23; 
  wire  _T_24; 
  wire  _T_25; 
  wire  _T_26; 
  wire  _T_27; 
  wire [10:0] _T_28; 
  wire [10:0] _T_30; 
  wire [7:0] _T_31; 
  wire [10:0] _GEN_18; 
  wire [10:0] _T_33; 
  wire  _T_41; 
  wire [10:0] _T_42; 
  wire [10:0] _T_44; 
  wire [10:0] _GEN_20; 
  wire [10:0] _T_48; 
  wire  first; 
  wire [10:0] _T_56; 
  wire  formatValid; 
  reg [2:0] _T_59; 
  reg [31:0] _RAND_5;
  wire [2:0] _GEN_7; 
  wire [7:0] formatOH; 
  wire  _T_60; 
  wire  _T_61; 
  wire  _T_62; 
  wire  _T_63; 
  wire  _T_64; 
  wire  _T_65; 
  wire  _T_69; 
  wire  _T_70; 
  wire  _T_72; 
  wire  _T_73; 
  wire  _T_75; 
  wire  _T_76; 
  wire  _T_78; 
  wire  _T_79; 
  wire  _T_81; 
  wire  _T_82; 
  wire  _T_84; 
  wire  _T_85; 
  wire  _T_87; 
  wire  _T_88; 
  wire  _T_90; 
  wire  _T_91; 
  wire  _T_93; 
  wire  _T_94; 
  wire  _T_96; 
  wire  _T_97; 
  reg [19:0] tx_a; 
  reg [31:0] _RAND_6;
  reg [19:0] tx_b; 
  reg [31:0] _RAND_7;
  reg [19:0] tx_c; 
  reg [31:0] _RAND_8;
  reg [19:0] tx_d; 
  reg [31:0] _RAND_9;
  reg [19:0] tx_e; 
  reg [31:0] _RAND_10;
  reg [19:0] rx_a; 
  reg [31:0] _RAND_11;
  reg [19:0] rx_b; 
  reg [31:0] _RAND_12;
  reg [19:0] rx_c; 
  reg [31:0] _RAND_13;
  reg [19:0] rx_d; 
  reg [31:0] _RAND_14;
  reg [19:0] rx_e; 
  reg [31:0] _RAND_15;
  wire  _T_100; 
  wire  _T_101; 
  wire  _T_102; 
  wire  _T_103; 
  wire  _T_104; 
  wire  _T_106; 
  wire [4:0] _T_108; 
  wire  _T_109; 
  wire [31:0] _T_112; 
  wire [20:0] _T_113; 
  wire [19:0] _T_114; 
  wire [19:0] _T_115; 
  wire [4:0] _T_116; 
  wire  _T_117; 
  wire [31:0] _T_120; 
  wire [20:0] _T_121; 
  wire [19:0] _T_122; 
  wire [19:0] _T_123; 
  wire [4:0] _T_124; 
  wire  _T_125; 
  wire [31:0] _T_128; 
  wire [20:0] _T_129; 
  wire [19:0] _T_130; 
  wire [19:0] _T_131; 
  wire [4:0] _T_132; 
  wire  _T_133; 
  wire [31:0] _T_136; 
  wire [20:0] _T_137; 
  wire [19:0] _T_138; 
  wire [19:0] _T_139; 
  wire [4:0] _T_140; 
  wire  _T_141; 
  wire [31:0] _T_144; 
  wire [20:0] _T_145; 
  wire [19:0] _T_146; 
  wire [19:0] _T_147; 
  wire [19:0] txInc_a; 
  wire [19:0] txInc_b; 
  wire [19:0] txInc_c; 
  wire [19:0] txInc_d; 
  wire [19:0] txInc_e; 
  wire [20:0] _T_150; 
  wire  _T_151; 
  wire [20:0] _T_154; 
  wire [20:0] _T_155; 
  wire  _T_156; 
  wire [20:0] _T_159; 
  wire [20:0] _T_160; 
  wire  _T_161; 
  wire [20:0] _T_164; 
  wire [20:0] _T_165; 
  wire  _T_166; 
  wire [20:0] _T_169; 
  wire [20:0] _T_170; 
  wire  _T_171; 
  wire [20:0] _T_174; 
  wire [19:0] rxInc_a; 
  wire [20:0] _T_176; 
  wire  _T_177; 
  wire [20:0] _T_180; 
  wire [19:0] rxInc_b; 
  wire [20:0] _T_181; 
  wire  _T_182; 
  wire [20:0] _T_185; 
  wire [19:0] rxInc_c; 
  wire [20:0] _T_186; 
  wire  _T_187; 
  wire [20:0] _T_190; 
  wire [19:0] rxInc_d; 
  wire [20:0] _T_191; 
  wire  _T_192; 
  wire [20:0] _T_195; 
  wire [19:0] rxInc_e; 
  wire [20:0] _T_196; 
  wire  _T_197; 
  wire [20:0] _T_200; 
  wire  txOut_ready; 
  wire [19:0] _T_149_a; 
  wire [19:0] _T_149_b; 
  wire [19:0] _T_149_c; 
  wire [19:0] _T_149_d; 
  wire [19:0] _T_149_e; 
  wire  rxOut_ready; 
  wire [19:0] _T_175_a; 
  wire [19:0] _T_175_b; 
  wire [19:0] _T_175_c; 
  wire [19:0] _T_175_d; 
  wire [19:0] _T_175_e; 
  dual_HellaQueue hqa ( 
    .clock(hqa_clock),
    .reset(hqa_reset),
    .io_enq_ready(hqa_io_enq_ready),
    .io_enq_valid(hqa_io_enq_valid),
    .io_enq_bits(hqa_io_enq_bits),
    .io_deq_ready(hqa_io_deq_ready),
    .io_deq_valid(hqa_io_deq_valid),
    .io_deq_bits(hqa_io_deq_bits)
  );
  dual_HellaQueue hqb ( 
    .clock(hqb_clock),
    .reset(hqb_reset),
    .io_enq_ready(hqb_io_enq_ready),
    .io_enq_valid(hqb_io_enq_valid),
    .io_enq_bits(hqb_io_enq_bits),
    .io_deq_ready(hqb_io_deq_ready),
    .io_deq_valid(hqb_io_deq_valid),
    .io_deq_bits(hqb_io_deq_bits)
  );
  dual_HellaQueue hqc ( 
    .clock(hqc_clock),
    .reset(hqc_reset),
    .io_enq_ready(hqc_io_enq_ready),
    .io_enq_valid(hqc_io_enq_valid),
    .io_enq_bits(hqc_io_enq_bits),
    .io_deq_ready(hqc_io_deq_ready),
    .io_deq_valid(hqc_io_deq_valid),
    .io_deq_bits(hqc_io_deq_bits)
  );
  dual_HellaQueue hqd ( 
    .clock(hqd_clock),
    .reset(hqd_reset),
    .io_enq_ready(hqd_io_enq_ready),
    .io_enq_valid(hqd_io_enq_valid),
    .io_enq_bits(hqd_io_enq_bits),
    .io_deq_ready(hqd_io_deq_ready),
    .io_deq_valid(hqd_io_deq_valid),
    .io_deq_bits(hqd_io_deq_bits)
  );
  dual_HellaQueue hqe ( 
    .clock(hqe_clock),
    .reset(hqe_reset),
    .io_enq_ready(hqe_io_enq_ready),
    .io_enq_valid(hqe_io_enq_valid),
    .io_enq_bits(hqe_io_enq_bits),
    .io_deq_ready(hqe_io_deq_ready),
    .io_deq_valid(hqe_io_deq_valid),
    .io_deq_bits(hqe_io_deq_bits)
  );
  dual_AsyncQueueSource AsyncQueueSource ( 
    .clock(AsyncQueueSource_clock),
    .reset(AsyncQueueSource_reset),
    .io_enq_ready(AsyncQueueSource_io_enq_ready),
    .io_enq_valid(AsyncQueueSource_io_enq_valid),
    .io_enq_bits(AsyncQueueSource_io_enq_bits),
    .io_async_mem_0(AsyncQueueSource_io_async_mem_0),
    .io_async_mem_1(AsyncQueueSource_io_async_mem_1),
    .io_async_mem_2(AsyncQueueSource_io_async_mem_2),
    .io_async_mem_3(AsyncQueueSource_io_async_mem_3),
    .io_async_mem_4(AsyncQueueSource_io_async_mem_4),
    .io_async_mem_5(AsyncQueueSource_io_async_mem_5),
    .io_async_mem_6(AsyncQueueSource_io_async_mem_6),
    .io_async_mem_7(AsyncQueueSource_io_async_mem_7),
    .io_async_ridx(AsyncQueueSource_io_async_ridx),
    .io_async_widx(AsyncQueueSource_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSource_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSource_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSource_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSource_io_async_safe_sink_reset_n)
  );
  dual_AsyncQueueSource AsyncQueueSource_1 ( 
    .clock(AsyncQueueSource_1_clock),
    .reset(AsyncQueueSource_1_reset),
    .io_enq_ready(AsyncQueueSource_1_io_enq_ready),
    .io_enq_valid(AsyncQueueSource_1_io_enq_valid),
    .io_enq_bits(AsyncQueueSource_1_io_enq_bits),
    .io_async_mem_0(AsyncQueueSource_1_io_async_mem_0),
    .io_async_mem_1(AsyncQueueSource_1_io_async_mem_1),
    .io_async_mem_2(AsyncQueueSource_1_io_async_mem_2),
    .io_async_mem_3(AsyncQueueSource_1_io_async_mem_3),
    .io_async_mem_4(AsyncQueueSource_1_io_async_mem_4),
    .io_async_mem_5(AsyncQueueSource_1_io_async_mem_5),
    .io_async_mem_6(AsyncQueueSource_1_io_async_mem_6),
    .io_async_mem_7(AsyncQueueSource_1_io_async_mem_7),
    .io_async_ridx(AsyncQueueSource_1_io_async_ridx),
    .io_async_widx(AsyncQueueSource_1_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSource_1_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSource_1_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSource_1_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSource_1_io_async_safe_sink_reset_n)
  );
  dual_AsyncQueueSource AsyncQueueSource_2 ( 
    .clock(AsyncQueueSource_2_clock),
    .reset(AsyncQueueSource_2_reset),
    .io_enq_ready(AsyncQueueSource_2_io_enq_ready),
    .io_enq_valid(AsyncQueueSource_2_io_enq_valid),
    .io_enq_bits(AsyncQueueSource_2_io_enq_bits),
    .io_async_mem_0(AsyncQueueSource_2_io_async_mem_0),
    .io_async_mem_1(AsyncQueueSource_2_io_async_mem_1),
    .io_async_mem_2(AsyncQueueSource_2_io_async_mem_2),
    .io_async_mem_3(AsyncQueueSource_2_io_async_mem_3),
    .io_async_mem_4(AsyncQueueSource_2_io_async_mem_4),
    .io_async_mem_5(AsyncQueueSource_2_io_async_mem_5),
    .io_async_mem_6(AsyncQueueSource_2_io_async_mem_6),
    .io_async_mem_7(AsyncQueueSource_2_io_async_mem_7),
    .io_async_ridx(AsyncQueueSource_2_io_async_ridx),
    .io_async_widx(AsyncQueueSource_2_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSource_2_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSource_2_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSource_2_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSource_2_io_async_safe_sink_reset_n)
  );
  dual_AsyncQueueSource AsyncQueueSource_3 ( 
    .clock(AsyncQueueSource_3_clock),
    .reset(AsyncQueueSource_3_reset),
    .io_enq_ready(AsyncQueueSource_3_io_enq_ready),
    .io_enq_valid(AsyncQueueSource_3_io_enq_valid),
    .io_enq_bits(AsyncQueueSource_3_io_enq_bits),
    .io_async_mem_0(AsyncQueueSource_3_io_async_mem_0),
    .io_async_mem_1(AsyncQueueSource_3_io_async_mem_1),
    .io_async_mem_2(AsyncQueueSource_3_io_async_mem_2),
    .io_async_mem_3(AsyncQueueSource_3_io_async_mem_3),
    .io_async_mem_4(AsyncQueueSource_3_io_async_mem_4),
    .io_async_mem_5(AsyncQueueSource_3_io_async_mem_5),
    .io_async_mem_6(AsyncQueueSource_3_io_async_mem_6),
    .io_async_mem_7(AsyncQueueSource_3_io_async_mem_7),
    .io_async_ridx(AsyncQueueSource_3_io_async_ridx),
    .io_async_widx(AsyncQueueSource_3_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSource_3_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSource_3_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSource_3_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSource_3_io_async_safe_sink_reset_n)
  );
  dual_AsyncQueueSource AsyncQueueSource_4 ( 
    .clock(AsyncQueueSource_4_clock),
    .reset(AsyncQueueSource_4_reset),
    .io_enq_ready(AsyncQueueSource_4_io_enq_ready),
    .io_enq_valid(AsyncQueueSource_4_io_enq_valid),
    .io_enq_bits(AsyncQueueSource_4_io_enq_bits),
    .io_async_mem_0(AsyncQueueSource_4_io_async_mem_0),
    .io_async_mem_1(AsyncQueueSource_4_io_async_mem_1),
    .io_async_mem_2(AsyncQueueSource_4_io_async_mem_2),
    .io_async_mem_3(AsyncQueueSource_4_io_async_mem_3),
    .io_async_mem_4(AsyncQueueSource_4_io_async_mem_4),
    .io_async_mem_5(AsyncQueueSource_4_io_async_mem_5),
    .io_async_mem_6(AsyncQueueSource_4_io_async_mem_6),
    .io_async_mem_7(AsyncQueueSource_4_io_async_mem_7),
    .io_async_ridx(AsyncQueueSource_4_io_async_ridx),
    .io_async_widx(AsyncQueueSource_4_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSource_4_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSource_4_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSource_4_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSource_4_io_async_safe_sink_reset_n)
  );
  dual_AsyncQueueSource_5 AsyncQueueSource_5 ( 
    .clock(AsyncQueueSource_5_clock),
    .reset(AsyncQueueSource_5_reset),
    .io_enq_ready(AsyncQueueSource_5_io_enq_ready),
    .io_enq_valid(AsyncQueueSource_5_io_enq_valid),
    .io_enq_bits_a(AsyncQueueSource_5_io_enq_bits_a),
    .io_enq_bits_b(AsyncQueueSource_5_io_enq_bits_b),
    .io_enq_bits_c(AsyncQueueSource_5_io_enq_bits_c),
    .io_enq_bits_d(AsyncQueueSource_5_io_enq_bits_d),
    .io_enq_bits_e(AsyncQueueSource_5_io_enq_bits_e),
    .io_async_mem_0_a(AsyncQueueSource_5_io_async_mem_0_a),
    .io_async_mem_0_b(AsyncQueueSource_5_io_async_mem_0_b),
    .io_async_mem_0_c(AsyncQueueSource_5_io_async_mem_0_c),
    .io_async_mem_0_d(AsyncQueueSource_5_io_async_mem_0_d),
    .io_async_mem_0_e(AsyncQueueSource_5_io_async_mem_0_e),
    .io_async_ridx(AsyncQueueSource_5_io_async_ridx),
    .io_async_widx(AsyncQueueSource_5_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSource_5_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSource_5_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSource_5_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSource_5_io_async_safe_sink_reset_n)
  );
  dual_AsyncQueueSource_5 AsyncQueueSource_6 ( 
    .clock(AsyncQueueSource_6_clock),
    .reset(AsyncQueueSource_6_reset),
    .io_enq_ready(AsyncQueueSource_6_io_enq_ready),
    .io_enq_valid(AsyncQueueSource_6_io_enq_valid),
    .io_enq_bits_a(AsyncQueueSource_6_io_enq_bits_a),
    .io_enq_bits_b(AsyncQueueSource_6_io_enq_bits_b),
    .io_enq_bits_c(AsyncQueueSource_6_io_enq_bits_c),
    .io_enq_bits_d(AsyncQueueSource_6_io_enq_bits_d),
    .io_enq_bits_e(AsyncQueueSource_6_io_enq_bits_e),
    .io_async_mem_0_a(AsyncQueueSource_6_io_async_mem_0_a),
    .io_async_mem_0_b(AsyncQueueSource_6_io_async_mem_0_b),
    .io_async_mem_0_c(AsyncQueueSource_6_io_async_mem_0_c),
    .io_async_mem_0_d(AsyncQueueSource_6_io_async_mem_0_d),
    .io_async_mem_0_e(AsyncQueueSource_6_io_async_mem_0_e),
    .io_async_ridx(AsyncQueueSource_6_io_async_ridx),
    .io_async_widx(AsyncQueueSource_6_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSource_6_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSource_6_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSource_6_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSource_6_io_async_safe_sink_reset_n)
  );
  assign _T_3 = b2c_data[2:0]; 
  assign _T_4 = b2c_data[5:3]; 
  assign _T_6 = b2c_data[12:9]; 
  assign _T_11 = 16'h1 << _T_6; 
  assign _T_12 = _T_11[12:0]; 
  assign _T_13 = _T_12[12:3]; 
  assign _T_14 = _T_6 <= 4'h2; 
  assign _T_15 = {_T_13,_T_14}; 
  assign _T_20 = _T_12[12:6]; 
  assign _T_21 = _T_6 <= 4'h5; 
  assign _T_22 = {_T_20,_T_21}; 
  assign _T_23 = _T_4 == 3'h4; 
  assign _T_24 = _T_4 == 3'h5; 
  assign _T_25 = _T_23 | _T_24; 
  assign _T_26 = _T_4 == 3'h1; 
  assign _T_27 = _T_4[2]; 
  assign _T_28 = _T_27 ? 11'h0 : _T_15; 
  assign _T_30 = _T_28 + 11'h2; 
  assign _T_31 = _T_26 ? _T_22 : 8'h0; 
  assign _GEN_18 = {{3'd0}, _T_31}; 
  assign _T_33 = _T_30 + _GEN_18; 
  assign _T_41 = _T_4[0]; 
  assign _T_42 = _T_41 ? _T_15 : 11'h0; 
  assign _T_44 = _T_42 + 11'h2; 
  assign _GEN_20 = {{10'd0}, _T_25}; 
  assign _T_48 = _T_42 + _GEN_20; 
  assign first = _T_2 == 11'h0; 
  assign _T_56 = _T_2 - 11'h1; 
  assign formatValid = b2c_send & first; 
  assign _GEN_7 = formatValid ? _T_3 : _T_59; 
  assign formatOH = 8'h1 << _GEN_7; 
  assign _T_60 = formatOH[0]; 
  assign _T_61 = formatOH[1]; 
  assign _T_62 = formatOH[2]; 
  assign _T_63 = formatOH[3]; 
  assign _T_64 = formatOH[4]; 
  assign _T_65 = formatOH[5]; 
  assign _T_69 = hqa_io_enq_valid == 1'h0; 
  assign _T_70 = _T_69 | hqa_io_enq_ready; 
  assign _T_72 = _T_70 | reset; 
  assign _T_73 = _T_72 == 1'h0; 
  assign _T_75 = hqb_io_enq_valid == 1'h0; 
  assign _T_76 = _T_75 | hqb_io_enq_ready; 
  assign _T_78 = _T_76 | reset; 
  assign _T_79 = _T_78 == 1'h0; 
  assign _T_81 = hqc_io_enq_valid == 1'h0; 
  assign _T_82 = _T_81 | hqc_io_enq_ready; 
  assign _T_84 = _T_82 | reset; 
  assign _T_85 = _T_84 == 1'h0; 
  assign _T_87 = hqd_io_enq_valid == 1'h0; 
  assign _T_88 = _T_87 | hqd_io_enq_ready; 
  assign _T_90 = _T_88 | reset; 
  assign _T_91 = _T_90 == 1'h0; 
  assign _T_93 = hqe_io_enq_valid == 1'h0; 
  assign _T_94 = _T_93 | hqe_io_enq_ready; 
  assign _T_96 = _T_94 | reset; 
  assign _T_97 = _T_96 == 1'h0; 
  assign _T_100 = hqa_io_deq_ready & hqa_io_deq_valid; 
  assign _T_101 = hqb_io_deq_ready & hqb_io_deq_valid; 
  assign _T_102 = hqc_io_deq_ready & hqc_io_deq_valid; 
  assign _T_103 = hqd_io_deq_ready & hqd_io_deq_valid; 
  assign _T_104 = hqe_io_deq_ready & hqe_io_deq_valid; 
  assign _T_106 = b2c_send & _T_65; 
  assign _T_108 = b2c_data[11:7]; 
  assign _T_109 = _T_108 > 5'h14; 
  assign _T_112 = 32'h1 << _T_108; 
  assign _T_113 = _T_112[20:0]; 
  assign _T_114 = _T_113[20:1]; 
  assign _T_115 = _T_109 ? 20'hfffff : _T_114; 
  assign _T_116 = b2c_data[16:12]; 
  assign _T_117 = _T_116 > 5'h14; 
  assign _T_120 = 32'h1 << _T_116; 
  assign _T_121 = _T_120[20:0]; 
  assign _T_122 = _T_121[20:1]; 
  assign _T_123 = _T_117 ? 20'hfffff : _T_122; 
  assign _T_124 = b2c_data[21:17]; 
  assign _T_125 = _T_124 > 5'h14; 
  assign _T_128 = 32'h1 << _T_124; 
  assign _T_129 = _T_128[20:0]; 
  assign _T_130 = _T_129[20:1]; 
  assign _T_131 = _T_125 ? 20'hfffff : _T_130; 
  assign _T_132 = b2c_data[26:22]; 
  assign _T_133 = _T_132 > 5'h14; 
  assign _T_136 = 32'h1 << _T_132; 
  assign _T_137 = _T_136[20:0]; 
  assign _T_138 = _T_137[20:1]; 
  assign _T_139 = _T_133 ? 20'hfffff : _T_138; 
  assign _T_140 = b2c_data[31:27]; 
  assign _T_141 = _T_140 > 5'h14; 
  assign _T_144 = 32'h1 << _T_140; 
  assign _T_145 = _T_144[20:0]; 
  assign _T_146 = _T_145[20:1]; 
  assign _T_147 = _T_141 ? 20'hfffff : _T_146; 
  assign txInc_a = _T_106 ? _T_115 : 20'h0; 
  assign txInc_b = _T_106 ? _T_123 : 20'h0; 
  assign txInc_c = _T_106 ? _T_131 : 20'h0; 
  assign txInc_d = _T_106 ? _T_139 : 20'h0; 
  assign txInc_e = _T_106 ? _T_147 : 20'h0; 
  assign _T_150 = tx_a + txInc_a; 
  assign _T_151 = _T_150[20:20]; 
  assign _T_154 = _T_151 ? 21'hfffff : _T_150; 
  assign _T_155 = tx_b + txInc_b; 
  assign _T_156 = _T_155[20:20]; 
  assign _T_159 = _T_156 ? 21'hfffff : _T_155; 
  assign _T_160 = tx_c + txInc_c; 
  assign _T_161 = _T_160[20:20]; 
  assign _T_164 = _T_161 ? 21'hfffff : _T_160; 
  assign _T_165 = tx_d + txInc_d; 
  assign _T_166 = _T_165[20:20]; 
  assign _T_169 = _T_166 ? 21'hfffff : _T_165; 
  assign _T_170 = tx_e + txInc_e; 
  assign _T_171 = _T_170[20:20]; 
  assign _T_174 = _T_171 ? 21'hfffff : _T_170; 
  assign rxInc_a = {{19'd0}, _T_100}; 
  assign _T_176 = rx_a + rxInc_a; 
  assign _T_177 = _T_176[20:20]; 
  assign _T_180 = _T_177 ? 21'hfffff : _T_176; 
  assign rxInc_b = {{19'd0}, _T_101}; 
  assign _T_181 = rx_b + rxInc_b; 
  assign _T_182 = _T_181[20:20]; 
  assign _T_185 = _T_182 ? 21'hfffff : _T_181; 
  assign rxInc_c = {{19'd0}, _T_102}; 
  assign _T_186 = rx_c + rxInc_c; 
  assign _T_187 = _T_186[20:20]; 
  assign _T_190 = _T_187 ? 21'hfffff : _T_186; 
  assign rxInc_d = {{19'd0}, _T_103}; 
  assign _T_191 = rx_d + rxInc_d; 
  assign _T_192 = _T_191[20:20]; 
  assign _T_195 = _T_192 ? 21'hfffff : _T_191; 
  assign rxInc_e = {{19'd0}, _T_104}; 
  assign _T_196 = rx_e + rxInc_e; 
  assign _T_197 = _T_196[20:20]; 
  assign _T_200 = _T_197 ? 21'hfffff : _T_196; 
  assign txOut_ready = AsyncQueueSource_5_io_enq_ready; 
  assign _T_149_a = _T_154[19:0]; 
  assign _T_149_b = _T_159[19:0]; 
  assign _T_149_c = _T_164[19:0]; 
  assign _T_149_d = _T_169[19:0]; 
  assign _T_149_e = _T_174[19:0]; 
  assign rxOut_ready = AsyncQueueSource_6_io_enq_ready; 
  assign _T_175_a = _T_180[19:0]; 
  assign _T_175_b = _T_185[19:0]; 
  assign _T_175_c = _T_190[19:0]; 
  assign _T_175_d = _T_195[19:0]; 
  assign _T_175_e = _T_200[19:0]; 
  assign io_a_mem_0 = AsyncQueueSource_io_async_mem_0; 
  assign io_a_mem_1 = AsyncQueueSource_io_async_mem_1; 
  assign io_a_mem_2 = AsyncQueueSource_io_async_mem_2; 
  assign io_a_mem_3 = AsyncQueueSource_io_async_mem_3; 
  assign io_a_mem_4 = AsyncQueueSource_io_async_mem_4; 
  assign io_a_mem_5 = AsyncQueueSource_io_async_mem_5; 
  assign io_a_mem_6 = AsyncQueueSource_io_async_mem_6; 
  assign io_a_mem_7 = AsyncQueueSource_io_async_mem_7; 
  assign io_a_widx = AsyncQueueSource_io_async_widx; 
  assign io_a_safe_widx_valid = AsyncQueueSource_io_async_safe_widx_valid; 
  assign io_a_safe_source_reset_n = AsyncQueueSource_io_async_safe_source_reset_n; 
  assign io_bmem_0 = AsyncQueueSource_1_io_async_mem_0; 
  assign io_bmem_1 = AsyncQueueSource_1_io_async_mem_1; 
  assign io_bmem_2 = AsyncQueueSource_1_io_async_mem_2; 
  assign io_bmem_3 = AsyncQueueSource_1_io_async_mem_3; 
  assign io_bmem_4 = AsyncQueueSource_1_io_async_mem_4; 
  assign io_bmem_5 = AsyncQueueSource_1_io_async_mem_5; 
  assign io_bmem_6 = AsyncQueueSource_1_io_async_mem_6; 
  assign io_bmem_7 = AsyncQueueSource_1_io_async_mem_7; 
  assign io_bwidx = AsyncQueueSource_1_io_async_widx; 
  assign io_bsafe_widx_valid = AsyncQueueSource_1_io_async_safe_widx_valid; 
  assign io_bsafe_source_reset_n = AsyncQueueSource_1_io_async_safe_source_reset_n; 
  assign io_c_mem_0 = AsyncQueueSource_2_io_async_mem_0; 
  assign io_c_mem_1 = AsyncQueueSource_2_io_async_mem_1; 
  assign io_c_mem_2 = AsyncQueueSource_2_io_async_mem_2; 
  assign io_c_mem_3 = AsyncQueueSource_2_io_async_mem_3; 
  assign io_c_mem_4 = AsyncQueueSource_2_io_async_mem_4; 
  assign io_c_mem_5 = AsyncQueueSource_2_io_async_mem_5; 
  assign io_c_mem_6 = AsyncQueueSource_2_io_async_mem_6; 
  assign io_c_mem_7 = AsyncQueueSource_2_io_async_mem_7; 
  assign io_c_widx = AsyncQueueSource_2_io_async_widx; 
  assign io_c_safe_widx_valid = AsyncQueueSource_2_io_async_safe_widx_valid; 
  assign io_c_safe_source_reset_n = AsyncQueueSource_2_io_async_safe_source_reset_n; 
  assign io_d_mem_0 = AsyncQueueSource_3_io_async_mem_0; 
  assign io_d_mem_1 = AsyncQueueSource_3_io_async_mem_1; 
  assign io_d_mem_2 = AsyncQueueSource_3_io_async_mem_2; 
  assign io_d_mem_3 = AsyncQueueSource_3_io_async_mem_3; 
  assign io_d_mem_4 = AsyncQueueSource_3_io_async_mem_4; 
  assign io_d_mem_5 = AsyncQueueSource_3_io_async_mem_5; 
  assign io_d_mem_6 = AsyncQueueSource_3_io_async_mem_6; 
  assign io_d_mem_7 = AsyncQueueSource_3_io_async_mem_7; 
  assign io_d_widx = AsyncQueueSource_3_io_async_widx; 
  assign io_d_safe_widx_valid = AsyncQueueSource_3_io_async_safe_widx_valid; 
  assign io_d_safe_source_reset_n = AsyncQueueSource_3_io_async_safe_source_reset_n; 
  assign io_e_mem_0 = AsyncQueueSource_4_io_async_mem_0; 
  assign io_e_mem_1 = AsyncQueueSource_4_io_async_mem_1; 
  assign io_e_mem_2 = AsyncQueueSource_4_io_async_mem_2; 
  assign io_e_mem_3 = AsyncQueueSource_4_io_async_mem_3; 
  assign io_e_mem_4 = AsyncQueueSource_4_io_async_mem_4; 
  assign io_e_mem_5 = AsyncQueueSource_4_io_async_mem_5; 
  assign io_e_mem_6 = AsyncQueueSource_4_io_async_mem_6; 
  assign io_e_mem_7 = AsyncQueueSource_4_io_async_mem_7; 
  assign io_e_widx = AsyncQueueSource_4_io_async_widx; 
  assign io_e_safe_widx_valid = AsyncQueueSource_4_io_async_safe_widx_valid; 
  assign io_e_safe_source_reset_n = AsyncQueueSource_4_io_async_safe_source_reset_n; 
  assign io_rxc_mem_0_a = AsyncQueueSource_6_io_async_mem_0_a; 
  assign io_rxc_mem_0_b = AsyncQueueSource_6_io_async_mem_0_b; 
  assign io_rxc_mem_0_c = AsyncQueueSource_6_io_async_mem_0_c; 
  assign io_rxc_mem_0_d = AsyncQueueSource_6_io_async_mem_0_d; 
  assign io_rxc_mem_0_e = AsyncQueueSource_6_io_async_mem_0_e; 
  assign io_rxc_widx = AsyncQueueSource_6_io_async_widx; 
  assign io_rxc_safe_widx_valid = AsyncQueueSource_6_io_async_safe_widx_valid; 
  assign io_rxc_safe_source_reset_n = AsyncQueueSource_6_io_async_safe_source_reset_n; 
  assign io_txc_mem_0_a = AsyncQueueSource_5_io_async_mem_0_a; 
  assign io_txc_mem_0_b = AsyncQueueSource_5_io_async_mem_0_b; 
  assign io_txc_mem_0_c = AsyncQueueSource_5_io_async_mem_0_c; 
  assign io_txc_mem_0_d = AsyncQueueSource_5_io_async_mem_0_d; 
  assign io_txc_mem_0_e = AsyncQueueSource_5_io_async_mem_0_e; 
  assign io_txc_widx = AsyncQueueSource_5_io_async_widx; 
  assign io_txc_safe_widx_valid = AsyncQueueSource_5_io_async_safe_widx_valid; 
  assign io_txc_safe_source_reset_n = AsyncQueueSource_5_io_async_safe_source_reset_n; 
  assign hqa_clock = clock; 
  assign hqa_reset = reset; 
  assign hqa_io_enq_valid = b2c_send & _T_60; 
  assign hqa_io_enq_bits = b2c_data; 
  assign hqa_io_deq_ready = AsyncQueueSource_io_enq_ready; 
  assign hqb_clock = clock; 
  assign hqb_reset = reset; 
  assign hqb_io_enq_valid = b2c_send & _T_61; 
  assign hqb_io_enq_bits = b2c_data; 
  assign hqb_io_deq_ready = AsyncQueueSource_1_io_enq_ready; 
  assign hqc_clock = clock; 
  assign hqc_reset = reset; 
  assign hqc_io_enq_valid = b2c_send & _T_62; 
  assign hqc_io_enq_bits = b2c_data; 
  assign hqc_io_deq_ready = AsyncQueueSource_2_io_enq_ready; 
  assign hqd_clock = clock; 
  assign hqd_reset = reset; 
  assign hqd_io_enq_valid = b2c_send & _T_63; 
  assign hqd_io_enq_bits = b2c_data; 
  assign hqd_io_deq_ready = AsyncQueueSource_3_io_enq_ready; 
  assign hqe_clock = clock; 
  assign hqe_reset = reset; 
  assign hqe_io_enq_valid = b2c_send & _T_64; 
  assign hqe_io_enq_bits = b2c_data; 
  assign hqe_io_deq_ready = AsyncQueueSource_4_io_enq_ready; 
  assign AsyncQueueSource_clock = clock; 
  assign AsyncQueueSource_reset = reset; 
  assign AsyncQueueSource_io_enq_valid = hqa_io_deq_valid; 
  assign AsyncQueueSource_io_enq_bits = hqa_io_deq_bits; 
  assign AsyncQueueSource_io_async_ridx = io_a_ridx; 
  assign AsyncQueueSource_io_async_safe_ridx_valid = io_a_safe_ridx_valid; 
  assign AsyncQueueSource_io_async_safe_sink_reset_n = io_a_safe_sink_reset_n; 
  assign AsyncQueueSource_1_clock = clock; 
  assign AsyncQueueSource_1_reset = reset; 
  assign AsyncQueueSource_1_io_enq_valid = hqb_io_deq_valid; 
  assign AsyncQueueSource_1_io_enq_bits = hqb_io_deq_bits; 
  assign AsyncQueueSource_1_io_async_ridx = io_bridx; 
  assign AsyncQueueSource_1_io_async_safe_ridx_valid = io_bsafe_ridx_valid; 
  assign AsyncQueueSource_1_io_async_safe_sink_reset_n = io_bsafe_sink_reset_n; 
  assign AsyncQueueSource_2_clock = clock; 
  assign AsyncQueueSource_2_reset = reset; 
  assign AsyncQueueSource_2_io_enq_valid = hqc_io_deq_valid; 
  assign AsyncQueueSource_2_io_enq_bits = hqc_io_deq_bits; 
  assign AsyncQueueSource_2_io_async_ridx = io_c_ridx; 
  assign AsyncQueueSource_2_io_async_safe_ridx_valid = io_c_safe_ridx_valid; 
  assign AsyncQueueSource_2_io_async_safe_sink_reset_n = io_c_safe_sink_reset_n; 
  assign AsyncQueueSource_3_clock = clock; 
  assign AsyncQueueSource_3_reset = reset; 
  assign AsyncQueueSource_3_io_enq_valid = hqd_io_deq_valid; 
  assign AsyncQueueSource_3_io_enq_bits = hqd_io_deq_bits; 
  assign AsyncQueueSource_3_io_async_ridx = io_d_ridx; 
  assign AsyncQueueSource_3_io_async_safe_ridx_valid = io_d_safe_ridx_valid; 
  assign AsyncQueueSource_3_io_async_safe_sink_reset_n = io_d_safe_sink_reset_n; 
  assign AsyncQueueSource_4_clock = clock; 
  assign AsyncQueueSource_4_reset = reset; 
  assign AsyncQueueSource_4_io_enq_valid = hqe_io_deq_valid; 
  assign AsyncQueueSource_4_io_enq_bits = hqe_io_deq_bits; 
  assign AsyncQueueSource_4_io_async_ridx = io_e_ridx; 
  assign AsyncQueueSource_4_io_async_safe_ridx_valid = io_e_safe_ridx_valid; 
  assign AsyncQueueSource_4_io_async_safe_sink_reset_n = io_e_safe_sink_reset_n; 
  assign AsyncQueueSource_5_clock = clock; 
  assign AsyncQueueSource_5_reset = reset; 
  assign AsyncQueueSource_5_io_enq_valid = 1'h1; 
  assign AsyncQueueSource_5_io_enq_bits_a = tx_a; 
  assign AsyncQueueSource_5_io_enq_bits_b = tx_b; 
  assign AsyncQueueSource_5_io_enq_bits_c = tx_c; 
  assign AsyncQueueSource_5_io_enq_bits_d = tx_d; 
  assign AsyncQueueSource_5_io_enq_bits_e = tx_e; 
  assign AsyncQueueSource_5_io_async_ridx = io_txc_ridx; 
  assign AsyncQueueSource_5_io_async_safe_ridx_valid = io_txc_safe_ridx_valid; 
  assign AsyncQueueSource_5_io_async_safe_sink_reset_n = io_txc_safe_sink_reset_n; 
  assign AsyncQueueSource_6_clock = clock; 
  assign AsyncQueueSource_6_reset = reset; 
  assign AsyncQueueSource_6_io_enq_valid = 1'h1; 
  assign AsyncQueueSource_6_io_enq_bits_a = rx_a; 
  assign AsyncQueueSource_6_io_enq_bits_b = rx_b; 
  assign AsyncQueueSource_6_io_enq_bits_c = rx_c; 
  assign AsyncQueueSource_6_io_enq_bits_d = rx_d; 
  assign AsyncQueueSource_6_io_enq_bits_e = rx_e; 
  assign AsyncQueueSource_6_io_async_ridx = io_rxc_ridx; 
  assign AsyncQueueSource_6_io_async_safe_ridx_valid = io_rxc_safe_ridx_valid; 
  assign AsyncQueueSource_6_io_async_safe_sink_reset_n = io_rxc_safe_sink_reset_n; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  b2c_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  b2c_send = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_2 = _RAND_4[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_59 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  tx_a = _RAND_6[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  tx_b = _RAND_7[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  tx_c = _RAND_8[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  tx_d = _RAND_9[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  tx_e = _RAND_10[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  rx_a = _RAND_11[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  rx_b = _RAND_12[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  rx_c = _RAND_13[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  rx_d = _RAND_14[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  rx_e = _RAND_15[19:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    _T <= io_b2c_data;
    b2c_data <= _T;
    _T_1 <= io_b2c_send;
    if (reset) begin
      b2c_send <= 1'h0;
    end else begin
      b2c_send <= _T_1;
    end
    if (reset) begin
      _T_2 <= 11'h0;
    end else begin
      if (b2c_send) begin
        if (first) begin
          if (3'h5 == _T_3) begin
            _T_2 <= 11'h0;
          end else begin
            if (3'h4 == _T_3) begin
              _T_2 <= 11'h0;
            end else begin
              if (3'h3 == _T_3) begin
                _T_2 <= _T_48;
              end else begin
                if (3'h2 == _T_3) begin
                  _T_2 <= _T_44;
                end else begin
                  if (3'h1 == _T_3) begin
                    _T_2 <= _T_33;
                  end else begin
                    _T_2 <= _T_33;
                  end
                end
              end
            end
          end
        end else begin
          _T_2 <= _T_56;
        end
      end
    end
    if (formatValid) begin
      _T_59 <= _T_3;
    end
    if (reset) begin
      tx_a <= 20'h0;
    end else begin
      if (txOut_ready) begin
        if (_T_106) begin
          if (_T_109) begin
            tx_a <= 20'hfffff;
          end else begin
            tx_a <= _T_114;
          end
        end else begin
          tx_a <= 20'h0;
        end
      end else begin
        tx_a <= _T_149_a;
      end
    end
    if (reset) begin
      tx_b <= 20'h0;
    end else begin
      if (txOut_ready) begin
        if (_T_106) begin
          if (_T_117) begin
            tx_b <= 20'hfffff;
          end else begin
            tx_b <= _T_122;
          end
        end else begin
          tx_b <= 20'h0;
        end
      end else begin
        tx_b <= _T_149_b;
      end
    end
    if (reset) begin
      tx_c <= 20'h0;
    end else begin
      if (txOut_ready) begin
        if (_T_106) begin
          if (_T_125) begin
            tx_c <= 20'hfffff;
          end else begin
            tx_c <= _T_130;
          end
        end else begin
          tx_c <= 20'h0;
        end
      end else begin
        tx_c <= _T_149_c;
      end
    end
    if (reset) begin
      tx_d <= 20'h0;
    end else begin
      if (txOut_ready) begin
        if (_T_106) begin
          if (_T_133) begin
            tx_d <= 20'hfffff;
          end else begin
            tx_d <= _T_138;
          end
        end else begin
          tx_d <= 20'h0;
        end
      end else begin
        tx_d <= _T_149_d;
      end
    end
    if (reset) begin
      tx_e <= 20'h0;
    end else begin
      if (txOut_ready) begin
        if (_T_106) begin
          if (_T_141) begin
            tx_e <= 20'hfffff;
          end else begin
            tx_e <= _T_146;
          end
        end else begin
          tx_e <= 20'h0;
        end
      end else begin
        tx_e <= _T_149_e;
      end
    end
    if (reset) begin
      rx_a <= 20'h800;
    end else begin
      if (rxOut_ready) begin
        rx_a <= rxInc_a;
      end else begin
        rx_a <= _T_175_a;
      end
    end
    if (reset) begin
      rx_b <= 20'h800;
    end else begin
      if (rxOut_ready) begin
        rx_b <= rxInc_b;
      end else begin
        rx_b <= _T_175_b;
      end
    end
    if (reset) begin
      rx_c <= 20'h800;
    end else begin
      if (rxOut_ready) begin
        rx_c <= rxInc_c;
      end else begin
        rx_c <= _T_175_c;
      end
    end
    if (reset) begin
      rx_d <= 20'h800;
    end else begin
      if (rxOut_ready) begin
        rx_d <= rxInc_d;
      end else begin
        rx_d <= _T_175_d;
      end
    end
    if (reset) begin
      rx_e <= 20'h800;
    end else begin
      if (rxOut_ready) begin
        rx_e <= rxInc_e;
      end else begin
        rx_e <= _T_175_e;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_73) begin
          $fwrite(32'h80000002,"Assertion failed\n    at dual_RX.scala:55 assert (!hq.io.enq.valid || hq.io.enq.ready) // overrun impossible\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_73) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_79) begin
          $fwrite(32'h80000002,"Assertion failed\n    at dual_RX.scala:55 assert (!hq.io.enq.valid || hq.io.enq.ready) // overrun impossible\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_79) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_85) begin
          $fwrite(32'h80000002,"Assertion failed\n    at dual_RX.scala:55 assert (!hq.io.enq.valid || hq.io.enq.ready) // overrun impossible\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_85) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_91) begin
          $fwrite(32'h80000002,"Assertion failed\n    at dual_RX.scala:55 assert (!hq.io.enq.valid || hq.io.enq.ready) // overrun impossible\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_91) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_97) begin
          $fwrite(32'h80000002,"Assertion failed\n    at dual_RX.scala:55 assert (!hq.io.enq.valid || hq.io.enq.ready) // overrun impossible\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_97) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_ShiftQueue( 
  input         clock, 
  input         reset, 
  output        io_enq_ready, 
  input         io_enq_valid, 
  input  [31:0] io_enq_bits_data, 
  input         io_enq_bits_last, 
  input  [12:0] io_enq_bits_beats, 
  input         io_deq_ready, 
  output        io_deq_valid, 
  output [31:0] io_deq_bits_data, 
  output        io_deq_bits_last, 
  output [12:0] io_deq_bits_beats 
);
  reg  _T_1_0; 
  reg [31:0] _RAND_0;
  reg  _T_1_1; 
  reg [31:0] _RAND_1;
  reg [31:0] _T_2_0_data; 
  reg [31:0] _RAND_2;
  reg  _T_2_0_last; 
  reg [31:0] _RAND_3;
  reg [12:0] _T_2_0_beats; 
  reg [31:0] _RAND_4;
  reg [31:0] _T_2_1_data; 
  reg [31:0] _RAND_5;
  reg  _T_2_1_last; 
  reg [31:0] _RAND_6;
  reg [12:0] _T_2_1_beats; 
  reg [31:0] _RAND_7;
  wire  _T_4; 
  wire  _T_7; 
  wire  _T_10; 
  wire  _T_11; 
  wire  _T_12; 
  wire  _T_19; 
  wire  _T_23; 
  wire  _T_26; 
  wire  _T_27; 
  wire  _T_28; 
  wire  _T_29; 
  wire  _T_36; 
  assign _T_4 = io_enq_ready & io_enq_valid; 
  assign _T_7 = _T_1_1 | _T_4; 
  assign _T_10 = _T_1_0 == 1'h0; 
  assign _T_11 = _T_4 & _T_10; 
  assign _T_12 = io_deq_ready ? _T_7 : _T_11; 
  assign _T_19 = _T_4 | _T_1_0; 
  assign _T_23 = _T_4 & _T_1_1; 
  assign _T_26 = _T_4 & _T_1_0; 
  assign _T_27 = _T_1_1 == 1'h0; 
  assign _T_28 = _T_26 & _T_27; 
  assign _T_29 = io_deq_ready ? _T_23 : _T_28; 
  assign _T_36 = _T_26 | _T_1_1; 
  assign io_enq_ready = _T_1_1 == 1'h0; 
  assign io_deq_valid = _T_1_0; 
  assign io_deq_bits_data = _T_2_0_data; 
  assign io_deq_bits_last = _T_2_0_last; 
  assign io_deq_bits_beats = _T_2_0_beats; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2_0_data = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_2_0_last = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_2_0_beats = _RAND_4[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_2_1_data = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_2_1_last = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_2_1_beats = _RAND_7[12:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_1_0 <= 1'h0;
    end else begin
      if (io_deq_ready) begin
        _T_1_0 <= _T_7;
      end else begin
        _T_1_0 <= _T_19;
      end
    end
    if (reset) begin
      _T_1_1 <= 1'h0;
    end else begin
      if (io_deq_ready) begin
        _T_1_1 <= _T_23;
      end else begin
        _T_1_1 <= _T_36;
      end
    end
    if (_T_12) begin
      if (_T_1_1) begin
        _T_2_0_data <= _T_2_1_data;
      end else begin
        _T_2_0_data <= io_enq_bits_data;
      end
    end
    if (_T_12) begin
      if (_T_1_1) begin
        _T_2_0_last <= _T_2_1_last;
      end else begin
        _T_2_0_last <= io_enq_bits_last;
      end
    end
    if (_T_12) begin
      if (_T_1_1) begin
        _T_2_0_beats <= _T_2_1_beats;
      end else begin
        _T_2_0_beats <= io_enq_bits_beats;
      end
    end
    if (_T_29) begin
      _T_2_1_data <= io_enq_bits_data;
    end
    if (_T_29) begin
      _T_2_1_last <= io_enq_bits_last;
    end
    if (_T_29) begin
      _T_2_1_beats <= io_enq_bits_beats;
    end
  end
endmodule
module dual_SinkA( 
  input         clock, 
  input         reset, 
  output        io_a_ready, 
  input         io_a_valid, 
  input  [2:0]  io_a_bits_opcode, 
  input  [2:0]  io_a_bits_param, 
  input  [2:0]  io_a_bits_size, 
  input  [2:0]  io_a_bits_source, 
  input  [31:0] io_a_bits_address, 
  input  [3:0]  io_a_bits_mask, 
  input  [31:0] io_a_bits_data, 
  input         io_q_ready, 
  output        io_q_valid, 
  output [31:0] io_q_bits_data, 
  output        io_q_bits_last, 
  output [12:0] io_q_bits_beats 
);
  wire  inject_clock; 
  wire  inject_reset; 
  wire  inject_io_i_last; 
  wire  inject_io_o_last; 
  wire  inject_io_i_ready; 
  wire  inject_io_i_valid; 
  wire [2:0] inject_io_i_bits_opcode; 
  wire [2:0] inject_io_i_bits_param; 
  wire [2:0] inject_io_i_bits_size; 
  wire [2:0] inject_io_i_bits_source; 
  wire [31:0] inject_io_i_bits_address; 
  wire [3:0] inject_io_i_bits_mask; 
  wire [31:0] inject_io_i_bits_data; 
  wire  inject_io_o_ready; 
  wire  inject_io_o_valid; 
  wire [2:0] inject_io_o_bits_opcode; 
  wire [2:0] inject_io_o_bits_param; 
  wire [2:0] inject_io_o_bits_size; 
  wire [2:0] inject_io_o_bits_source; 
  wire [31:0] inject_io_o_bits_address; 
  wire [31:0] inject_io_o_bits_data; 
  wire  Queue_clock; 
  wire  Queue_reset; 
  wire  Queue_io_enq_ready; 
  wire  Queue_io_enq_valid; 
  wire [2:0] Queue_io_enq_bits_opcode; 
  wire [2:0] Queue_io_enq_bits_param; 
  wire [2:0] Queue_io_enq_bits_size; 
  wire [2:0] Queue_io_enq_bits_source; 
  wire [31:0] Queue_io_enq_bits_address; 
  wire [3:0] Queue_io_enq_bits_mask; 
  wire [31:0] Queue_io_enq_bits_data; 
  wire  Queue_io_deq_ready; 
  wire  Queue_io_deq_valid; 
  wire [2:0] Queue_io_deq_bits_opcode; 
  wire [2:0] Queue_io_deq_bits_param; 
  wire [2:0] Queue_io_deq_bits_size; 
  wire [2:0] Queue_io_deq_bits_source; 
  wire [31:0] Queue_io_deq_bits_address; 
  wire [3:0] Queue_io_deq_bits_mask; 
  wire [31:0] Queue_io_deq_bits_data; 
  wire  _T; 
  wire [12:0] _T_2; 
  wire [5:0] _T_3; 
  wire [5:0] _T_4; 
  wire [3:0] _T_5; 
  wire  _T_6; 
  wire  _T_7; 
  wire [3:0] _T_8; 
  reg [3:0] _T_9; 
  reg [31:0] _RAND_0;
  wire [3:0] _T_11; 
  wire  _T_12; 
  wire  _T_13; 
  wire  _T_14; 
  wire  _T_20; 
  wire  a_hasData; 
  wire  a_partial; 
  reg [1:0] state; 
  reg [31:0] _RAND_1;
  wire  _T_21; 
  wire  _T_22; 
  wire  _T_23; 
  wire  _T_24; 
  wire  _T_26; 
  wire  _T_27; 
  wire [1:0] _GEN_7; 
  wire [1:0] _GEN_8; 
  wire [1:0] _GEN_9; 
  wire [1:0] _GEN_10; 
  wire [1:0] _GEN_11; 
  wire [1:0] _GEN_12; 
  wire [1:0] _GEN_13; 
  wire [15:0] _T_29; 
  wire [1:0] _GEN_18; 
  wire [1:0] _GEN_19; 
  wire [1:0] _GEN_20; 
  wire [1:0] _GEN_21; 
  wire [2:0] _T_31; 
  wire [3:0] _T_33; 
  wire [2:0] _T_35; 
  wire [2:0] _T_37; 
  wire [31:0] header; 
  wire [1:0] _T_45; 
  wire  isLastState; 
  wire [31:0] _T_48_1; 
  wire [31:0] _GEN_23; 
  wire [31:0] _GEN_24; 
  wire [31:0] _T_48_3; 
  wire [15:0] _T_51; 
  wire [12:0] _T_52; 
  wire [9:0] _T_53; 
  wire  _T_54; 
  wire [10:0] _T_55; 
  wire [10:0] _T_56; 
  wire [10:0] _T_58; 
  wire [6:0] _T_63; 
  wire  _T_64; 
  wire [7:0] _T_65; 
  wire [7:0] _T_66; 
  wire [10:0] _GEN_26; 
  wire [10:0] _T_68; 
  dual_PartialInjector inject ( 
    .clock(inject_clock),
    .reset(inject_reset),
    .io_i_last(inject_io_i_last),
    .io_o_last(inject_io_o_last),
    .io_i_ready(inject_io_i_ready),
    .io_i_valid(inject_io_i_valid),
    .io_i_bits_opcode(inject_io_i_bits_opcode),
    .io_i_bits_param(inject_io_i_bits_param),
    .io_i_bits_size(inject_io_i_bits_size),
    .io_i_bits_source(inject_io_i_bits_source),
    .io_i_bits_address(inject_io_i_bits_address),
    .io_i_bits_mask(inject_io_i_bits_mask),
    .io_i_bits_data(inject_io_i_bits_data),
    .io_o_ready(inject_io_o_ready),
    .io_o_valid(inject_io_o_valid),
    .io_o_bits_opcode(inject_io_o_bits_opcode),
    .io_o_bits_param(inject_io_o_bits_param),
    .io_o_bits_size(inject_io_o_bits_size),
    .io_o_bits_source(inject_io_o_bits_source),
    .io_o_bits_address(inject_io_o_bits_address),
    .io_o_bits_data(inject_io_o_bits_data)
  );
  dual_Queue_5 dual_Queue ( 
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_opcode(Queue_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_io_enq_bits_param),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_source(Queue_io_enq_bits_source),
    .io_enq_bits_address(Queue_io_enq_bits_address),
    .io_enq_bits_mask(Queue_io_enq_bits_mask),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_opcode(Queue_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_io_deq_bits_param),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_source(Queue_io_deq_bits_source),
    .io_deq_bits_address(Queue_io_deq_bits_address),
    .io_deq_bits_mask(Queue_io_deq_bits_mask),
    .io_deq_bits_data(Queue_io_deq_bits_data)
  );
  assign _T = inject_io_i_ready & inject_io_i_valid; 
  assign _T_2 = 13'h3f << inject_io_i_bits_size; 
  assign _T_3 = _T_2[5:0]; 
  assign _T_4 = ~ _T_3; 
  assign _T_5 = _T_4[5:2]; 
  assign _T_6 = inject_io_i_bits_opcode[2]; 
  assign _T_7 = _T_6 == 1'h0; 
  assign _T_8 = _T_7 ? _T_5 : 4'h0; 
  assign _T_11 = _T_9 - 4'h1; 
  assign _T_12 = _T_9 == 4'h0; 
  assign _T_13 = _T_9 == 4'h1; 
  assign _T_14 = _T_8 == 4'h0; 
  assign _T_20 = inject_io_o_bits_opcode[2]; 
  assign a_hasData = _T_20 == 1'h0; 
  assign a_partial = inject_io_o_bits_opcode == 3'h1; 
  assign _T_21 = io_q_ready & io_q_valid; 
  assign _T_22 = 2'h0 == state; 
  assign _T_23 = 2'h1 == state; 
  assign _T_24 = 2'h2 == state; 
  assign _T_26 = 2'h3 == state; 
  assign _T_27 = inject_io_o_last == 1'h0; 
  assign _GEN_7 = 3'h1 == inject_io_o_bits_source ? 2'h1 : 2'h0; 
  assign _GEN_8 = 3'h2 == inject_io_o_bits_source ? 2'h2 : _GEN_7; 
  assign _GEN_9 = 3'h3 == inject_io_o_bits_source ? 2'h3 : _GEN_8; 
  assign _GEN_10 = 3'h4 == inject_io_o_bits_source ? 2'h0 : _GEN_9; 
  assign _GEN_11 = 3'h5 == inject_io_o_bits_source ? 2'h1 : _GEN_10; 
  assign _GEN_12 = 3'h6 == inject_io_o_bits_source ? 2'h2 : _GEN_11; 
  assign _GEN_13 = 3'h7 == inject_io_o_bits_source ? 2'h3 : _GEN_12; 
  assign _T_29 = {{14'd0}, _GEN_13}; 
  assign _GEN_18 = 3'h4 == inject_io_o_bits_source ? 2'h2 : 2'h1; 
  assign _GEN_19 = 3'h5 == inject_io_o_bits_source ? 2'h2 : _GEN_18; 
  assign _GEN_20 = 3'h6 == inject_io_o_bits_source ? 2'h2 : _GEN_19; 
  assign _GEN_21 = 3'h7 == inject_io_o_bits_source ? 2'h2 : _GEN_20; 
  assign _T_31 = {{1'd0}, _GEN_21}; 
  assign _T_33 = {{1'd0}, inject_io_o_bits_size}; 
  assign _T_35 = inject_io_o_bits_param; 
  assign _T_37 = inject_io_o_bits_opcode; 
  assign header = {_T_29,_T_31,_T_33,_T_35,_T_37,3'h0}; 
  assign _T_45 = a_hasData ? 2'h3 : 2'h2; 
  assign isLastState = state == _T_45; 
  assign _T_48_1 = inject_io_o_bits_address; 
  assign _GEN_23 = 2'h1 == state ? _T_48_1 : header; 
  assign _GEN_24 = 2'h2 == state ? 32'h0 : _GEN_23; 
  assign _T_48_3 = inject_io_o_bits_data; 
  assign _T_51 = 16'h1 << _T_33; 
  assign _T_52 = _T_51[12:0]; 
  assign _T_53 = _T_52[12:3]; 
  assign _T_54 = inject_io_o_bits_size <= 3'h2; 
  assign _T_55 = {_T_53,_T_54}; 
  assign _T_56 = a_hasData ? _T_55 : 11'h0; 
  assign _T_58 = _T_56 + 11'h3; 
  assign _T_63 = _T_52[12:6]; 
  assign _T_64 = inject_io_o_bits_size <= 3'h5; 
  assign _T_65 = {_T_63,_T_64}; 
  assign _T_66 = a_partial ? _T_65 : 8'h0; 
  assign _GEN_26 = {{3'd0}, _T_66}; 
  assign _T_68 = _T_58 + _GEN_26; 
  assign io_a_ready = Queue_io_enq_ready; 
  assign io_q_valid = inject_io_o_valid; 
  assign io_q_bits_data = 2'h3 == state ? _T_48_3 : _GEN_24; 
  assign io_q_bits_last = inject_io_o_last & isLastState; 
  assign io_q_bits_beats = {{2'd0}, _T_68}; 
  assign inject_clock = clock; 
  assign inject_reset = reset; 
  assign inject_io_i_last = _T_13 | _T_14; 
  assign inject_io_i_valid = Queue_io_deq_valid; 
  assign inject_io_i_bits_opcode = Queue_io_deq_bits_opcode; 
  assign inject_io_i_bits_param = Queue_io_deq_bits_param; 
  assign inject_io_i_bits_size = Queue_io_deq_bits_size; 
  assign inject_io_i_bits_source = Queue_io_deq_bits_source; 
  assign inject_io_i_bits_address = Queue_io_deq_bits_address; 
  assign inject_io_i_bits_mask = Queue_io_deq_bits_mask; 
  assign inject_io_i_bits_data = Queue_io_deq_bits_data; 
  assign inject_io_o_ready = io_q_ready & isLastState; 
  assign Queue_clock = clock; 
  assign Queue_reset = reset; 
  assign Queue_io_enq_valid = io_a_valid; 
  assign Queue_io_enq_bits_opcode = io_a_bits_opcode; 
  assign Queue_io_enq_bits_param = io_a_bits_param; 
  assign Queue_io_enq_bits_size = io_a_bits_size; 
  assign Queue_io_enq_bits_source = io_a_bits_source; 
  assign Queue_io_enq_bits_address = io_a_bits_address; 
  assign Queue_io_enq_bits_mask = io_a_bits_mask; 
  assign Queue_io_enq_bits_data = io_a_bits_data; 
  assign Queue_io_deq_ready = inject_io_i_ready; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_9 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_9 <= 4'h0;
    end else begin
      if (_T) begin
        if (_T_12) begin
          if (_T_7) begin
            _T_9 <= _T_5;
          end else begin
            _T_9 <= 4'h0;
          end
        end else begin
          _T_9 <= _T_11;
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_21) begin
        if (_T_22) begin
          state <= 2'h1;
        end else begin
          if (_T_23) begin
            state <= 2'h2;
          end else begin
            if (_T_24) begin
              if (a_hasData) begin
                state <= 2'h3;
              end else begin
                state <= 2'h0;
              end
            end else begin
              if (_T_26) begin
                if (_T_27) begin
                  state <= 2'h3;
                end else begin
                  state <= 2'h0;
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module dual_SinkB( 
  input         clock, 
  input         reset, 
  input         io_q_ready, 
  output        io_q_valid, 
  output [31:0] io_q_bits_data, 
  output        io_q_bits_last 
);
  reg [1:0] state; 
  reg [31:0] _RAND_0;
  wire  _T_22; 
  wire  _T_23; 
  wire  _T_24; 
  wire  _T_25; 
  wire  _T_27; 
  wire [31:0] _GEN_7; 
  wire [31:0] _GEN_8; 
  assign _T_22 = io_q_ready & io_q_valid; 
  assign _T_23 = 2'h0 == state; 
  assign _T_24 = 2'h1 == state; 
  assign _T_25 = 2'h2 == state; 
  assign _T_27 = 2'h3 == state; 
  assign _GEN_7 = 2'h1 == state ? 32'h0 : 32'h1; 
  assign _GEN_8 = 2'h2 == state ? 32'h0 : _GEN_7; 
  assign io_q_valid = 1'h0; 
  assign io_q_bits_data = 2'h3 == state ? 32'h0 : _GEN_8; 
  assign io_q_bits_last = state == 2'h2; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_22) begin
        if (_T_23) begin
          state <= 2'h1;
        end else begin
          if (_T_24) begin
            state <= 2'h2;
          end else begin
            if (_T_25) begin
              state <= 2'h0;
            end else begin
              if (_T_27) begin
                state <= 2'h0;
              end
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at dual_SinkB.scala:48 assert (!b.valid || b.bits.source === UInt(0))\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_SinkC( 
  input         clock, 
  input         reset, 
  input         io_q_ready, 
  output        io_q_valid, 
  output [31:0] io_q_bits_data, 
  output        io_q_bits_last 
);
  reg [1:0] state; 
  reg [31:0] _RAND_0;
  wire  _T_21; 
  wire  _T_22; 
  wire  _T_23; 
  wire  _T_24; 
  wire  _T_26; 
  wire [31:0] _GEN_23; 
  wire [31:0] _GEN_24; 
  assign _T_21 = io_q_ready & io_q_valid; 
  assign _T_22 = 2'h0 == state; 
  assign _T_23 = 2'h1 == state; 
  assign _T_24 = 2'h2 == state; 
  assign _T_26 = 2'h3 == state; 
  assign _GEN_23 = 2'h1 == state ? 32'h0 : 32'h2; 
  assign _GEN_24 = 2'h2 == state ? 32'h0 : _GEN_23; 
  assign io_q_valid = 1'h0; 
  assign io_q_bits_data = 2'h3 == state ? 32'h0 : _GEN_24; 
  assign io_q_bits_last = state == 2'h2; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_21) begin
        if (_T_22) begin
          state <= 2'h1;
        end else begin
          if (_T_23) begin
            state <= 2'h2;
          end else begin
            if (_T_24) begin
              state <= 2'h0;
            end else begin
              if (_T_26) begin
                state <= 2'h0;
              end
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at dual_SinkC.scala:50 assert (!c.valid || domain(c.bits.source) === UInt(0))\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_SinkD( 
  input         clock, 
  input         reset, 
  output        io_d_ready, 
  input         io_d_valid, 
  input  [2:0]  io_d_bits_opcode, 
  input  [1:0]  io_d_bits_param, 
  input  [3:0]  io_d_bits_size, 
  input  [5:0]  io_d_bits_source, 
  input         io_d_bits_sink, 
  input         io_d_bits_denied, 
  input  [31:0] io_d_bits_data, 
  input         io_q_ready, 
  output        io_q_valid, 
  output [31:0] io_q_bits_data, 
  output        io_q_bits_last, 
  output [12:0] io_q_bits_beats, 
  output        io_a_tlSource_valid, 
  output [5:0]  io_a_tlSource_bits, 
  input  [15:0] io_a_clSource, 
  output        io_c_tlSource_valid, 
  output [5:0]  io_c_tlSource_bits, 
  input  [15:0] io_c_clSource 
);
  wire  d_clock; 
  wire  d_reset; 
  wire  d_io_enq_ready; 
  wire  d_io_enq_valid; 
  wire [2:0] d_io_enq_bits_opcode; 
  wire [1:0] d_io_enq_bits_param; 
  wire [3:0] d_io_enq_bits_size; 
  wire [5:0] d_io_enq_bits_source; 
  wire  d_io_enq_bits_sink; 
  wire  d_io_enq_bits_denied; 
  wire [31:0] d_io_enq_bits_data; 
  wire  d_io_deq_ready; 
  wire  d_io_deq_valid; 
  wire [2:0] d_io_deq_bits_opcode; 
  wire [1:0] d_io_deq_bits_param; 
  wire [3:0] d_io_deq_bits_size; 
  wire [5:0] d_io_deq_bits_source; 
  wire  d_io_deq_bits_sink; 
  wire  d_io_deq_bits_denied; 
  wire [31:0] d_io_deq_bits_data; 
  reg [1:0] state; 
  reg [31:0] _RAND_0;
  wire  _T; 
  wire [22:0] _T_2; 
  wire [7:0] _T_3; 
  wire [7:0] _T_4; 
  wire [5:0] _T_5; 
  wire  _T_6; 
  wire [5:0] _T_7; 
  reg [5:0] _T_8; 
  reg [31:0] _RAND_1;
  wire [5:0] _T_10; 
  wire  _T_11; 
  wire  _T_12; 
  wire  _T_13; 
  wire  d_last; 
  wire  _T_18; 
  wire  _T_19; 
  wire  d_grant; 
  wire  _T_20; 
  wire  _T_21; 
  wire  _T_24; 
  wire  _T_26; 
  wire  relack; 
  wire  _T_29; 
  wire  _T_30; 
  wire  _T_31; 
  wire [2:0] _T_38; 
  wire [15:0] _T_39; 
  wire [3:0] _T_44; 
  wire [2:0] _T_48; 
  wire [31:0] header; 
  wire [1:0] _T_56; 
  wire [1:0] _T_57; 
  wire  isLastState; 
  wire [31:0] _T_60_1; 
  wire [31:0] _GEN_6; 
  wire [31:0] _T_60_2; 
  wire [15:0] _T_63; 
  wire [12:0] _T_64; 
  wire [9:0] _T_65; 
  wire  _T_66; 
  wire [10:0] _T_67; 
  wire [10:0] _T_68; 
  wire [10:0] _T_70; 
  wire [10:0] _GEN_8; 
  wire [10:0] _T_72; 
  dual_Queue_8 d ( 
    .clock(d_clock),
    .reset(d_reset),
    .io_enq_ready(d_io_enq_ready),
    .io_enq_valid(d_io_enq_valid),
    .io_enq_bits_opcode(d_io_enq_bits_opcode),
    .io_enq_bits_param(d_io_enq_bits_param),
    .io_enq_bits_size(d_io_enq_bits_size),
    .io_enq_bits_source(d_io_enq_bits_source),
    .io_enq_bits_sink(d_io_enq_bits_sink),
    .io_enq_bits_denied(d_io_enq_bits_denied),
    .io_enq_bits_data(d_io_enq_bits_data),
    .io_deq_ready(d_io_deq_ready),
    .io_deq_valid(d_io_deq_valid),
    .io_deq_bits_opcode(d_io_deq_bits_opcode),
    .io_deq_bits_param(d_io_deq_bits_param),
    .io_deq_bits_size(d_io_deq_bits_size),
    .io_deq_bits_source(d_io_deq_bits_source),
    .io_deq_bits_sink(d_io_deq_bits_sink),
    .io_deq_bits_denied(d_io_deq_bits_denied),
    .io_deq_bits_data(d_io_deq_bits_data)
  );
  assign _T = d_io_deq_ready & d_io_deq_valid; 
  assign _T_2 = 23'hff << d_io_deq_bits_size; 
  assign _T_3 = _T_2[7:0]; 
  assign _T_4 = ~ _T_3; 
  assign _T_5 = _T_4[7:2]; 
  assign _T_6 = d_io_deq_bits_opcode[0]; 
  assign _T_7 = _T_6 ? _T_5 : 6'h0; 
  assign _T_10 = _T_8 - 6'h1; 
  assign _T_11 = _T_8 == 6'h0; 
  assign _T_12 = _T_8 == 6'h1; 
  assign _T_13 = _T_7 == 6'h0; 
  assign d_last = _T_12 | _T_13; 
  assign _T_18 = d_io_deq_bits_opcode == 3'h4; 
  assign _T_19 = d_io_deq_bits_opcode == 3'h5; 
  assign d_grant = _T_18 | _T_19; 
  assign _T_20 = io_q_ready & io_q_valid; 
  assign _T_21 = 2'h0 == state; 
  assign _T_24 = 2'h1 == state; 
  assign _T_26 = 2'h2 == state; 
  assign relack = d_io_deq_bits_opcode == 3'h6; 
  assign _T_29 = state == 2'h0; 
  assign _T_30 = _T_20 & _T_29; 
  assign _T_31 = relack == 1'h0; 
  assign _T_38 = d_io_deq_bits_source[5:3]; 
  assign _T_39 = relack ? io_c_clSource : io_a_clSource; 
  assign _T_44 = d_io_deq_bits_size; 
  assign _T_48 = d_io_deq_bits_opcode; 
  assign header = {_T_39,_T_38,_T_44,d_io_deq_bits_denied,d_io_deq_bits_param,_T_48,3'h3}; 
  assign _T_56 = d_grant ? 2'h1 : 2'h0; 
  assign _T_57 = _T_6 ? 2'h2 : _T_56; 
  assign isLastState = state == _T_57; 
  assign _T_60_1 = {{31'd0}, d_io_deq_bits_sink}; 
  assign _GEN_6 = 2'h1 == state ? _T_60_1 : header; 
  assign _T_60_2 = d_io_deq_bits_data; 
  assign _T_63 = 16'h1 << _T_44; 
  assign _T_64 = _T_63[12:0]; 
  assign _T_65 = _T_64[12:3]; 
  assign _T_66 = d_io_deq_bits_size <= 4'h2; 
  assign _T_67 = {_T_65,_T_66}; 
  assign _T_68 = _T_6 ? _T_67 : 11'h0; 
  assign _T_70 = _T_68 + 11'h1; 
  assign _GEN_8 = {{10'd0}, d_grant}; 
  assign _T_72 = _T_70 + _GEN_8; 
  assign io_d_ready = d_io_enq_ready; 
  assign io_q_valid = d_io_deq_valid; 
  assign io_q_bits_data = 2'h2 == state ? _T_60_2 : _GEN_6; 
  assign io_q_bits_last = d_last & isLastState; 
  assign io_q_bits_beats = {{2'd0}, _T_72}; 
  assign io_a_tlSource_valid = _T_30 & _T_31; 
  assign io_a_tlSource_bits = d_io_deq_bits_source; 
  assign io_c_tlSource_valid = _T_30 & relack; 
  assign io_c_tlSource_bits = d_io_deq_bits_source; 
  assign d_clock = clock; 
  assign d_reset = reset; 
  assign d_io_enq_valid = io_d_valid; 
  assign d_io_enq_bits_opcode = io_d_bits_opcode; 
  assign d_io_enq_bits_param = io_d_bits_param; 
  assign d_io_enq_bits_size = io_d_bits_size; 
  assign d_io_enq_bits_source = io_d_bits_source; 
  assign d_io_enq_bits_sink = io_d_bits_sink; 
  assign d_io_enq_bits_denied = io_d_bits_denied; 
  assign d_io_enq_bits_data = io_d_bits_data; 
  assign d_io_deq_ready = io_q_ready & isLastState; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_8 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (d_grant) begin
            state <= 2'h1;
          end else begin
            if (_T_6) begin
              state <= 2'h2;
            end else begin
              state <= 2'h0;
            end
          end
        end else begin
          if (_T_24) begin
            if (_T_6) begin
              state <= 2'h2;
            end else begin
              state <= 2'h0;
            end
          end else begin
            if (_T_26) begin
              if (d_last) begin
                state <= 2'h0;
              end else begin
                state <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_8 <= 6'h0;
    end else begin
      if (_T) begin
        if (_T_11) begin
          if (_T_6) begin
            _T_8 <= _T_5;
          end else begin
            _T_8 <= 6'h0;
          end
        end else begin
          _T_8 <= _T_10;
        end
      end
    end
  end
endmodule
module dual_SinkE( 
  output [31:0] io_q_bits_data, 
  input  [15:0] io_d_clSink 
);
  wire [22:0] _T_16; 
  assign _T_16 = {io_d_clSink,3'h0,4'h0}; 
  assign io_q_bits_data = {_T_16,9'h4}; 
endmodule
module dual_SourceA( 
  input         clock, 
  input         reset, 
  input         io_a_ready, 
  output        io_a_valid, 
  output [2:0]  io_a_bits_opcode, 
  output [2:0]  io_a_bits_param, 
  output [3:0]  io_a_bits_size, 
  output [5:0]  io_a_bits_source, 
  output [31:0] io_a_bits_address, 
  output [3:0]  io_a_bits_mask, 
  output [31:0] io_a_bits_data, 
  output        io_q_ready, 
  input         io_q_valid, 
  input  [31:0] io_q_bits, 
  input         io_d_tlSource_valid, 
  input  [5:0]  io_d_tlSource_bits, 
  output [15:0] io_d_clSource 
);
  wire  cams_0_clock; 
  wire  cams_0_reset; 
  wire  cams_0_io_alloc_ready; 
  wire  cams_0_io_alloc_valid; 
  wire [15:0] cams_0_io_alloc_bits; 
  wire [2:0] cams_0_io_key; 
  wire  cams_0_io_free_valid; 
  wire [2:0] cams_0_io_free_bits; 
  wire [15:0] cams_0_io_data; 
  wire  cams_1_clock; 
  wire  cams_1_reset; 
  wire  cams_1_io_alloc_ready; 
  wire  cams_1_io_alloc_valid; 
  wire [15:0] cams_1_io_alloc_bits; 
  wire [2:0] cams_1_io_key; 
  wire  cams_1_io_free_valid; 
  wire [2:0] cams_1_io_free_bits; 
  wire [15:0] cams_1_io_data; 
  wire  cams_2_clock; 
  wire  cams_2_reset; 
  wire  cams_2_io_alloc_ready; 
  wire  cams_2_io_alloc_valid; 
  wire [15:0] cams_2_io_alloc_bits; 
  wire [2:0] cams_2_io_key; 
  wire  cams_2_io_free_valid; 
  wire [2:0] cams_2_io_free_bits; 
  wire [15:0] cams_2_io_data; 
  wire  cams_3_clock; 
  wire  cams_3_reset; 
  wire  cams_3_io_alloc_ready; 
  wire  cams_3_io_alloc_valid; 
  wire [15:0] cams_3_io_alloc_bits; 
  wire [2:0] cams_3_io_key; 
  wire  cams_3_io_free_valid; 
  wire [2:0] cams_3_io_free_bits; 
  wire [15:0] cams_3_io_data; 
  wire  cams_4_clock; 
  wire  cams_4_reset; 
  wire  cams_4_io_alloc_ready; 
  wire  cams_4_io_alloc_valid; 
  wire [15:0] cams_4_io_alloc_bits; 
  wire [2:0] cams_4_io_key; 
  wire  cams_4_io_free_valid; 
  wire [2:0] cams_4_io_free_bits; 
  wire [15:0] cams_4_io_data; 
  wire  cams_5_clock; 
  wire  cams_5_reset; 
  wire  cams_5_io_alloc_ready; 
  wire  cams_5_io_alloc_valid; 
  wire [15:0] cams_5_io_alloc_bits; 
  wire [2:0] cams_5_io_key; 
  wire  cams_5_io_free_valid; 
  wire [2:0] cams_5_io_free_bits; 
  wire [15:0] cams_5_io_data; 
  wire  cams_6_clock; 
  wire  cams_6_reset; 
  wire  cams_6_io_alloc_ready; 
  wire  cams_6_io_alloc_valid; 
  wire [15:0] cams_6_io_alloc_bits; 
  wire [2:0] cams_6_io_key; 
  wire  cams_6_io_free_valid; 
  wire [2:0] cams_6_io_free_bits; 
  wire [15:0] cams_6_io_data; 
  wire  cams_7_clock; 
  wire  cams_7_reset; 
  wire  cams_7_io_alloc_ready; 
  wire  cams_7_io_alloc_valid; 
  wire [15:0] cams_7_io_alloc_bits; 
  wire [2:0] cams_7_io_key; 
  wire  cams_7_io_free_valid; 
  wire [2:0] cams_7_io_free_bits; 
  wire [15:0] cams_7_io_data; 
  wire  extract_clock; 
  wire  extract_reset; 
  wire  extract_io_last; 
  wire  extract_io_i_ready; 
  wire  extract_io_i_valid; 
  wire [2:0] extract_io_i_bits_opcode; 
  wire [2:0] extract_io_i_bits_param; 
  wire [3:0] extract_io_i_bits_size; 
  wire [5:0] extract_io_i_bits_source; 
  wire [31:0] extract_io_i_bits_address; 
  wire [3:0] extract_io_i_bits_mask; 
  wire [31:0] extract_io_i_bits_data; 
  wire  extract_io_o_ready; 
  wire  extract_io_o_valid; 
  wire [2:0] extract_io_o_bits_opcode; 
  wire [2:0] extract_io_o_bits_param; 
  wire [3:0] extract_io_o_bits_size; 
  wire [5:0] extract_io_o_bits_source; 
  wire [31:0] extract_io_o_bits_address; 
  wire [3:0] extract_io_o_bits_mask; 
  wire [31:0] extract_io_o_bits_data; 
  reg [1:0] state; 
  reg [31:0] _RAND_0;
  wire [2:0] _T_1; 
  wire [2:0] _T_2; 
  wire [3:0] _T_3; 
  wire [2:0] _T_4; 
  wire [15:0] _T_5; 
  wire  _T_6; 
  reg [2:0] _T_10; 
  reg [31:0] _RAND_1;
  wire [2:0] _GEN_1; 
  reg [2:0] _T_12; 
  reg [31:0] _RAND_2;
  reg [3:0] _T_14; 
  reg [31:0] _RAND_3;
  wire [3:0] _GEN_3; 
  reg [2:0] _T_16; 
  reg [31:0] _RAND_4;
  wire [2:0] _GEN_4; 
  reg [15:0] _T_18; 
  reg [31:0] _RAND_5;
  wire  _T_19; 
  reg [31:0] _T_20; 
  reg [31:0] _RAND_6;
  wire [31:0] _GEN_6; 
  wire  _T_21; 
  reg [31:0] _T_22; 
  reg [31:0] _RAND_7;
  wire [31:0] _GEN_7; 
  reg [10:0] _T_23; 
  reg [31:0] _RAND_8;
  wire [15:0] _T_32; 
  wire [12:0] _T_33; 
  wire [9:0] _T_34; 
  wire  _T_35; 
  wire [10:0] _T_36; 
  wire [6:0] _T_41; 
  wire  _T_42; 
  wire [7:0] _T_43; 
  wire  _T_47; 
  wire  _T_48; 
  wire [10:0] _T_49; 
  wire [10:0] _T_51; 
  wire [7:0] _T_52; 
  wire [10:0] _GEN_40; 
  wire [10:0] _T_54; 
  wire  _T_71; 
  wire  _T_72; 
  wire  _T_73; 
  wire  _T_74; 
  wire  q_last; 
  wire  _T_75; 
  wire [10:0] _T_77; 
  wire  _T_79; 
  wire  q_hasData; 
  wire  _T_80; 
  reg  a_first; 
  reg [31:0] _RAND_9;
  wire  _T_83; 
  wire  _T_84; 
  wire  _T_85; 
  wire  _T_87; 
  wire  _T_88; 
  wire [63:0] q_address; 
  wire  _T_90; 
  wire  _T_91; 
  wire  q_acq; 
  wire [63:0] _T_95; 
  wire [64:0] _T_96; 
  wire [64:0] _T_97; 
  wire [64:0] _T_98; 
  wire  _T_99; 
  wire [63:0] _T_100; 
  wire [64:0] _T_101; 
  wire [64:0] _T_102; 
  wire [64:0] _T_103; 
  wire  _T_104; 
  wire [63:0] _T_105; 
  wire [64:0] _T_106; 
  wire [64:0] _T_107; 
  wire [64:0] _T_108; 
  wire  _T_109; 
  wire  _T_111; 
  wire  exists; 
  wire [64:0] _T_113; 
  wire [64:0] _T_130; 
  wire [64:0] _T_131; 
  wire  acquireOk; 
  wire  _T_139; 
  wire  _T_140; 
  wire  q_legal; 
  reg [2:0] _T_143; 
  reg [31:0] _RAND_10;
  wire [2:0] _T_142_0; 
  wire [2:0] _T_142_1; 
  wire [2:0] _GEN_16; 
  wire [2:0] _T_142_2; 
  wire [2:0] _GEN_17; 
  wire [2:0] _T_142_3; 
  wire [2:0] _GEN_18; 
  wire [2:0] _T_142_4; 
  wire [2:0] _GEN_19; 
  wire [2:0] _T_142_5; 
  wire [2:0] _GEN_20; 
  wire [2:0] _T_142_6; 
  wire [2:0] _GEN_21; 
  wire [2:0] _T_142_7; 
  wire [2:0] _GEN_22; 
  wire [2:0] _GEN_23; 
  wire [7:0] a_sel; 
  wire [63:0] _T_145; 
  wire [35:0] _T_146; 
  wire [27:0] _T_147; 
  wire [63:0] _T_148; 
  wire  _T_150; 
  wire [1:0] _T_151; 
  wire [1:0] _T_153; 
  wire  _T_154; 
  wire  _T_155; 
  wire  _T_156; 
  wire  _T_157; 
  wire  _T_159; 
  wire  _T_160; 
  wire  _T_162; 
  wire  _T_163; 
  wire  _T_164; 
  wire  _T_165; 
  wire  _T_166; 
  wire  _T_167; 
  wire  _T_168; 
  wire  _T_169; 
  wire  _T_170; 
  wire  _T_171; 
  wire  _T_172; 
  wire  _T_173; 
  wire  _T_174; 
  wire  _T_175; 
  wire  _T_176; 
  wire  _T_177; 
  wire  _T_178; 
  wire [1:0] _T_179; 
  wire [1:0] _T_180; 
  wire  _T_141_0; 
  wire  _T_141_1; 
  wire  _GEN_25; 
  wire  _T_141_2; 
  wire  _GEN_26; 
  wire  _T_141_3; 
  wire  _GEN_27; 
  wire  _T_141_4; 
  wire  _GEN_28; 
  wire  _T_141_5; 
  wire  _GEN_29; 
  wire  _T_141_6; 
  wire  _GEN_30; 
  wire  _T_141_7; 
  wire  _GEN_31; 
  wire  _T_182; 
  wire  stall; 
  wire  _T_183; 
  wire  xmit; 
  wire  _T_184; 
  wire  _T_185; 
  wire  _T_188; 
  wire  _T_189; 
  wire  _T_191; 
  wire  _T_192; 
  wire  _T_193; 
  wire  _T_194; 
  wire  _T_195; 
  wire  _T_196; 
  wire  _T_197; 
  wire  _T_198; 
  wire  _T_199; 
  wire  _T_200; 
  wire  _T_201; 
  wire  _T_203; 
  wire  _T_204; 
  wire  _T_205; 
  wire  _T_207; 
  wire  _T_208; 
  wire  _T_209; 
  wire  _T_211; 
  wire  _T_212; 
  wire  _T_213; 
  wire  _T_215; 
  wire  _T_216; 
  wire  _T_217; 
  wire  _T_219; 
  wire  _T_220; 
  wire  _T_221; 
  wire  _T_223; 
  wire  _T_224; 
  wire  _T_225; 
  wire  _T_227; 
  wire  _T_228; 
  wire  _T_229; 
  wire [2:0] d_clDomain; 
  wire [7:0] d_sel; 
  wire [15:0] _T_231_0; 
  wire [15:0] _T_231_1; 
  wire [15:0] _GEN_33; 
  wire [15:0] _T_231_2; 
  wire [15:0] _GEN_34; 
  wire [15:0] _T_231_3; 
  wire [15:0] _GEN_35; 
  wire [15:0] _T_231_4; 
  wire [15:0] _GEN_36; 
  wire [15:0] _T_231_5; 
  wire [15:0] _GEN_37; 
  wire [15:0] _T_231_6; 
  wire [15:0] _GEN_38; 
  wire [15:0] _T_231_7; 
  wire  _T_232; 
  wire  _T_233; 
  wire  _T_234; 
  wire  _T_235; 
  wire  _T_236; 
  wire  _T_237; 
  wire  _T_238; 
  wire  _T_239; 
  dual_CAM cams_0 ( 
    .clock(cams_0_clock),
    .reset(cams_0_reset),
    .io_alloc_ready(cams_0_io_alloc_ready),
    .io_alloc_valid(cams_0_io_alloc_valid),
    .io_alloc_bits(cams_0_io_alloc_bits),
    .io_key(cams_0_io_key),
    .io_free_valid(cams_0_io_free_valid),
    .io_free_bits(cams_0_io_free_bits),
    .io_data(cams_0_io_data)
  );
  dual_CAM cams_1 ( 
    .clock(cams_1_clock),
    .reset(cams_1_reset),
    .io_alloc_ready(cams_1_io_alloc_ready),
    .io_alloc_valid(cams_1_io_alloc_valid),
    .io_alloc_bits(cams_1_io_alloc_bits),
    .io_key(cams_1_io_key),
    .io_free_valid(cams_1_io_free_valid),
    .io_free_bits(cams_1_io_free_bits),
    .io_data(cams_1_io_data)
  );
  dual_CAM cams_2 ( 
    .clock(cams_2_clock),
    .reset(cams_2_reset),
    .io_alloc_ready(cams_2_io_alloc_ready),
    .io_alloc_valid(cams_2_io_alloc_valid),
    .io_alloc_bits(cams_2_io_alloc_bits),
    .io_key(cams_2_io_key),
    .io_free_valid(cams_2_io_free_valid),
    .io_free_bits(cams_2_io_free_bits),
    .io_data(cams_2_io_data)
  );
  dual_CAM cams_3 ( 
    .clock(cams_3_clock),
    .reset(cams_3_reset),
    .io_alloc_ready(cams_3_io_alloc_ready),
    .io_alloc_valid(cams_3_io_alloc_valid),
    .io_alloc_bits(cams_3_io_alloc_bits),
    .io_key(cams_3_io_key),
    .io_free_valid(cams_3_io_free_valid),
    .io_free_bits(cams_3_io_free_bits),
    .io_data(cams_3_io_data)
  );
  dual_CAM cams_4 ( 
    .clock(cams_4_clock),
    .reset(cams_4_reset),
    .io_alloc_ready(cams_4_io_alloc_ready),
    .io_alloc_valid(cams_4_io_alloc_valid),
    .io_alloc_bits(cams_4_io_alloc_bits),
    .io_key(cams_4_io_key),
    .io_free_valid(cams_4_io_free_valid),
    .io_free_bits(cams_4_io_free_bits),
    .io_data(cams_4_io_data)
  );
  dual_CAM cams_5 ( 
    .clock(cams_5_clock),
    .reset(cams_5_reset),
    .io_alloc_ready(cams_5_io_alloc_ready),
    .io_alloc_valid(cams_5_io_alloc_valid),
    .io_alloc_bits(cams_5_io_alloc_bits),
    .io_key(cams_5_io_key),
    .io_free_valid(cams_5_io_free_valid),
    .io_free_bits(cams_5_io_free_bits),
    .io_data(cams_5_io_data)
  );
  dual_CAM cams_6 ( 
    .clock(cams_6_clock),
    .reset(cams_6_reset),
    .io_alloc_ready(cams_6_io_alloc_ready),
    .io_alloc_valid(cams_6_io_alloc_valid),
    .io_alloc_bits(cams_6_io_alloc_bits),
    .io_key(cams_6_io_key),
    .io_free_valid(cams_6_io_free_valid),
    .io_free_bits(cams_6_io_free_bits),
    .io_data(cams_6_io_data)
  );
  dual_CAM cams_7 ( 
    .clock(cams_7_clock),
    .reset(cams_7_reset),
    .io_alloc_ready(cams_7_io_alloc_ready),
    .io_alloc_valid(cams_7_io_alloc_valid),
    .io_alloc_bits(cams_7_io_alloc_bits),
    .io_key(cams_7_io_key),
    .io_free_valid(cams_7_io_free_valid),
    .io_free_bits(cams_7_io_free_bits),
    .io_data(cams_7_io_data)
  );
  dual_ParitalExtractor extract ( 
    .clock(extract_clock),
    .reset(extract_reset),
    .io_last(extract_io_last),
    .io_i_ready(extract_io_i_ready),
    .io_i_valid(extract_io_i_valid),
    .io_i_bits_opcode(extract_io_i_bits_opcode),
    .io_i_bits_param(extract_io_i_bits_param),
    .io_i_bits_size(extract_io_i_bits_size),
    .io_i_bits_source(extract_io_i_bits_source),
    .io_i_bits_address(extract_io_i_bits_address),
    .io_i_bits_mask(extract_io_i_bits_mask),
    .io_i_bits_data(extract_io_i_bits_data),
    .io_o_ready(extract_io_o_ready),
    .io_o_valid(extract_io_o_valid),
    .io_o_bits_opcode(extract_io_o_bits_opcode),
    .io_o_bits_param(extract_io_o_bits_param),
    .io_o_bits_size(extract_io_o_bits_size),
    .io_o_bits_source(extract_io_o_bits_source),
    .io_o_bits_address(extract_io_o_bits_address),
    .io_o_bits_mask(extract_io_o_bits_mask),
    .io_o_bits_data(extract_io_o_bits_data)
  );
  assign _T_1 = io_q_bits[5:3]; 
  assign _T_2 = io_q_bits[8:6]; 
  assign _T_3 = io_q_bits[12:9]; 
  assign _T_4 = io_q_bits[15:13]; 
  assign _T_5 = io_q_bits[31:16]; 
  assign _T_6 = state == 2'h0; 
  assign _GEN_1 = _T_6 ? _T_1 : _T_10; 
  assign _GEN_3 = _T_6 ? _T_3 : _T_14; 
  assign _GEN_4 = _T_6 ? _T_4 : _T_16; 
  assign _T_19 = state == 2'h1; 
  assign _GEN_6 = _T_19 ? io_q_bits : _T_20; 
  assign _T_21 = state == 2'h2; 
  assign _GEN_7 = _T_21 ? io_q_bits : _T_22; 
  assign _T_32 = 16'h1 << _T_3; 
  assign _T_33 = _T_32[12:0]; 
  assign _T_34 = _T_33[12:3]; 
  assign _T_35 = _T_3 <= 4'h2; 
  assign _T_36 = {_T_34,_T_35}; 
  assign _T_41 = _T_33[12:6]; 
  assign _T_42 = _T_3 <= 4'h5; 
  assign _T_43 = {_T_41,_T_42}; 
  assign _T_47 = _T_1 == 3'h1; 
  assign _T_48 = _T_1[2]; 
  assign _T_49 = _T_48 ? 11'h0 : _T_36; 
  assign _T_51 = _T_49 + 11'h2; 
  assign _T_52 = _T_47 ? _T_43 : 8'h0; 
  assign _GEN_40 = {{3'd0}, _T_52}; 
  assign _T_54 = _T_51 + _GEN_40; 
  assign _T_71 = _T_23 == 11'h0; 
  assign _T_72 = _T_23 == 11'h1; 
  assign _T_73 = _T_54 == 11'h0; 
  assign _T_74 = _T_71 & _T_73; 
  assign q_last = _T_72 | _T_74; 
  assign _T_75 = io_q_ready & io_q_valid; 
  assign _T_77 = _T_23 - 11'h1; 
  assign _T_79 = _GEN_1[2]; 
  assign q_hasData = _T_79 == 1'h0; 
  assign _T_80 = state != 2'h3; 
  assign _T_83 = 2'h0 == state; 
  assign _T_84 = 2'h1 == state; 
  assign _T_85 = 2'h2 == state; 
  assign _T_87 = 2'h3 == state; 
  assign _T_88 = q_last == 1'h0; 
  assign q_address = {_GEN_7,_GEN_6}; 
  assign _T_90 = _GEN_1 == 3'h6; 
  assign _T_91 = _GEN_1 == 3'h7; 
  assign q_acq = _T_90 | _T_91; 
  assign _T_95 = q_address ^ 64'h80000000; 
  assign _T_96 = {1'b0,$signed(_T_95)}; 
  assign _T_97 = $signed(_T_96) & $signed(-65'sh80000000); 
  assign _T_98 = $signed(_T_97); 
  assign _T_99 = $signed(_T_98) == $signed(65'sh0); 
  assign _T_100 = q_address ^ 64'h40000000; 
  assign _T_101 = {1'b0,$signed(_T_100)}; 
  assign _T_102 = $signed(_T_101) & $signed(-65'sh20000000); 
  assign _T_103 = $signed(_T_102); 
  assign _T_104 = $signed(_T_103) == $signed(65'sh0); 
  assign _T_105 = q_address ^ 64'h10000000; 
  assign _T_106 = {1'b0,$signed(_T_105)}; 
  assign _T_107 = $signed(_T_106) & $signed(-65'sh10000000); 
  assign _T_108 = $signed(_T_107); 
  assign _T_109 = $signed(_T_108) == $signed(65'sh0); 
  assign _T_111 = _T_99 | _T_104; 
  assign exists = _T_111 | _T_109; 
  assign _T_113 = {1'b0,$signed(q_address)}; 
  assign _T_130 = $signed(_T_113) & $signed(65'shc0000000); 
  assign _T_131 = $signed(_T_130); 
  assign acquireOk = $signed(_T_131) == $signed(65'sh0); 
  assign _T_139 = q_acq == 1'h0; 
  assign _T_140 = _T_139 | acquireOk; 
  assign q_legal = exists & _T_140; 
  assign _T_142_0 = cams_0_io_key; 
  assign _T_142_1 = cams_1_io_key; 
  assign _GEN_16 = 3'h1 == _GEN_4 ? _T_142_1 : _T_142_0; 
  assign _T_142_2 = cams_2_io_key; 
  assign _GEN_17 = 3'h2 == _GEN_4 ? _T_142_2 : _GEN_16; 
  assign _T_142_3 = cams_3_io_key; 
  assign _GEN_18 = 3'h3 == _GEN_4 ? _T_142_3 : _GEN_17; 
  assign _T_142_4 = cams_4_io_key; 
  assign _GEN_19 = 3'h4 == _GEN_4 ? _T_142_4 : _GEN_18; 
  assign _T_142_5 = cams_5_io_key; 
  assign _GEN_20 = 3'h5 == _GEN_4 ? _T_142_5 : _GEN_19; 
  assign _T_142_6 = cams_6_io_key; 
  assign _GEN_21 = 3'h6 == _GEN_4 ? _T_142_6 : _GEN_20; 
  assign _T_142_7 = cams_7_io_key; 
  assign _GEN_22 = 3'h7 == _GEN_4 ? _T_142_7 : _GEN_21; 
  assign _GEN_23 = a_first ? _GEN_22 : _T_143; 
  assign a_sel = 8'h1 << _GEN_4; 
  assign _T_145 = q_legal ? q_address : 64'h10000000; 
  assign _T_146 = _T_145[63:28]; 
  assign _T_147 = q_address[27:0]; 
  assign _T_148 = {_T_146,_T_147}; 
  assign _T_150 = _GEN_3[0]; 
  assign _T_151 = 2'h1 << _T_150; 
  assign _T_153 = _T_151 | 2'h1; 
  assign _T_154 = _GEN_3 >= 4'h2; 
  assign _T_155 = _T_153[1]; 
  assign _T_156 = _GEN_6[1]; 
  assign _T_157 = _T_156 == 1'h0; 
  assign _T_159 = _T_155 & _T_157; 
  assign _T_160 = _T_154 | _T_159; 
  assign _T_162 = _T_155 & _T_156; 
  assign _T_163 = _T_154 | _T_162; 
  assign _T_164 = _T_153[0]; 
  assign _T_165 = _GEN_6[0]; 
  assign _T_166 = _T_165 == 1'h0; 
  assign _T_167 = _T_157 & _T_166; 
  assign _T_168 = _T_164 & _T_167; 
  assign _T_169 = _T_160 | _T_168; 
  assign _T_170 = _T_157 & _T_165; 
  assign _T_171 = _T_164 & _T_170; 
  assign _T_172 = _T_160 | _T_171; 
  assign _T_173 = _T_156 & _T_166; 
  assign _T_174 = _T_164 & _T_173; 
  assign _T_175 = _T_163 | _T_174; 
  assign _T_176 = _T_156 & _T_165; 
  assign _T_177 = _T_164 & _T_176; 
  assign _T_178 = _T_163 | _T_177; 
  assign _T_179 = {_T_172,_T_169}; 
  assign _T_180 = {_T_178,_T_175}; 
  assign _T_141_0 = cams_0_io_alloc_ready; 
  assign _T_141_1 = cams_1_io_alloc_ready; 
  assign _GEN_25 = 3'h1 == _GEN_4 ? _T_141_1 : _T_141_0; 
  assign _T_141_2 = cams_2_io_alloc_ready; 
  assign _GEN_26 = 3'h2 == _GEN_4 ? _T_141_2 : _GEN_25; 
  assign _T_141_3 = cams_3_io_alloc_ready; 
  assign _GEN_27 = 3'h3 == _GEN_4 ? _T_141_3 : _GEN_26; 
  assign _T_141_4 = cams_4_io_alloc_ready; 
  assign _GEN_28 = 3'h4 == _GEN_4 ? _T_141_4 : _GEN_27; 
  assign _T_141_5 = cams_5_io_alloc_ready; 
  assign _GEN_29 = 3'h5 == _GEN_4 ? _T_141_5 : _GEN_28; 
  assign _T_141_6 = cams_6_io_alloc_ready; 
  assign _GEN_30 = 3'h6 == _GEN_4 ? _T_141_6 : _GEN_29; 
  assign _T_141_7 = cams_7_io_alloc_ready; 
  assign _GEN_31 = 3'h7 == _GEN_4 ? _T_141_7 : _GEN_30; 
  assign _T_182 = _GEN_31 == 1'h0; 
  assign stall = a_first & _T_182; 
  assign _T_183 = state == 2'h3; 
  assign xmit = q_last | _T_183; 
  assign _T_184 = stall == 1'h0; 
  assign _T_185 = io_q_valid & _T_184; 
  assign _T_188 = extract_io_i_ready & _T_184; 
  assign _T_189 = xmit == 1'h0; 
  assign _T_191 = a_sel[0]; 
  assign _T_192 = a_sel[1]; 
  assign _T_193 = a_sel[2]; 
  assign _T_194 = a_sel[3]; 
  assign _T_195 = a_sel[4]; 
  assign _T_196 = a_sel[5]; 
  assign _T_197 = a_sel[6]; 
  assign _T_198 = a_sel[7]; 
  assign _T_199 = _T_191 & a_first; 
  assign _T_200 = _T_199 & xmit; 
  assign _T_201 = _T_200 & io_q_valid; 
  assign _T_203 = _T_192 & a_first; 
  assign _T_204 = _T_203 & xmit; 
  assign _T_205 = _T_204 & io_q_valid; 
  assign _T_207 = _T_193 & a_first; 
  assign _T_208 = _T_207 & xmit; 
  assign _T_209 = _T_208 & io_q_valid; 
  assign _T_211 = _T_194 & a_first; 
  assign _T_212 = _T_211 & xmit; 
  assign _T_213 = _T_212 & io_q_valid; 
  assign _T_215 = _T_195 & a_first; 
  assign _T_216 = _T_215 & xmit; 
  assign _T_217 = _T_216 & io_q_valid; 
  assign _T_219 = _T_196 & a_first; 
  assign _T_220 = _T_219 & xmit; 
  assign _T_221 = _T_220 & io_q_valid; 
  assign _T_223 = _T_197 & a_first; 
  assign _T_224 = _T_223 & xmit; 
  assign _T_225 = _T_224 & io_q_valid; 
  assign _T_227 = _T_198 & a_first; 
  assign _T_228 = _T_227 & xmit; 
  assign _T_229 = _T_228 & io_q_valid; 
  assign d_clDomain = io_d_tlSource_bits[5:3]; 
  assign d_sel = 8'h1 << d_clDomain; 
  assign _T_231_0 = cams_0_io_data; 
  assign _T_231_1 = cams_1_io_data; 
  assign _GEN_33 = 3'h1 == d_clDomain ? _T_231_1 : _T_231_0; 
  assign _T_231_2 = cams_2_io_data; 
  assign _GEN_34 = 3'h2 == d_clDomain ? _T_231_2 : _GEN_33; 
  assign _T_231_3 = cams_3_io_data; 
  assign _GEN_35 = 3'h3 == d_clDomain ? _T_231_3 : _GEN_34; 
  assign _T_231_4 = cams_4_io_data; 
  assign _GEN_36 = 3'h4 == d_clDomain ? _T_231_4 : _GEN_35; 
  assign _T_231_5 = cams_5_io_data; 
  assign _GEN_37 = 3'h5 == d_clDomain ? _T_231_5 : _GEN_36; 
  assign _T_231_6 = cams_6_io_data; 
  assign _GEN_38 = 3'h6 == d_clDomain ? _T_231_6 : _GEN_37; 
  assign _T_231_7 = cams_7_io_data; 
  assign _T_232 = d_sel[0]; 
  assign _T_233 = d_sel[1]; 
  assign _T_234 = d_sel[2]; 
  assign _T_235 = d_sel[3]; 
  assign _T_236 = d_sel[4]; 
  assign _T_237 = d_sel[5]; 
  assign _T_238 = d_sel[6]; 
  assign _T_239 = d_sel[7]; 
  assign io_a_valid = extract_io_o_valid; 
  assign io_a_bits_opcode = extract_io_o_bits_opcode; 
  assign io_a_bits_param = extract_io_o_bits_param; 
  assign io_a_bits_size = extract_io_o_bits_size; 
  assign io_a_bits_source = extract_io_o_bits_source; 
  assign io_a_bits_address = extract_io_o_bits_address; 
  assign io_a_bits_mask = extract_io_o_bits_mask; 
  assign io_a_bits_data = extract_io_o_bits_data; 
  assign io_q_ready = _T_188 | _T_189; 
  assign io_d_clSource = 3'h7 == d_clDomain ? _T_231_7 : _GEN_38; 
  assign cams_0_clock = clock; 
  assign cams_0_reset = reset; 
  assign cams_0_io_alloc_valid = _T_201 & extract_io_i_ready; 
  assign cams_0_io_alloc_bits = _T_6 ? _T_5 : _T_18; 
  assign cams_0_io_free_valid = io_d_tlSource_valid & _T_232; 
  assign cams_0_io_free_bits = io_d_tlSource_bits[2:0]; 
  assign cams_1_clock = clock; 
  assign cams_1_reset = reset; 
  assign cams_1_io_alloc_valid = _T_205 & extract_io_i_ready; 
  assign cams_1_io_alloc_bits = _T_6 ? _T_5 : _T_18; 
  assign cams_1_io_free_valid = io_d_tlSource_valid & _T_233; 
  assign cams_1_io_free_bits = io_d_tlSource_bits[2:0]; 
  assign cams_2_clock = clock; 
  assign cams_2_reset = reset; 
  assign cams_2_io_alloc_valid = _T_209 & extract_io_i_ready; 
  assign cams_2_io_alloc_bits = _T_6 ? _T_5 : _T_18; 
  assign cams_2_io_free_valid = io_d_tlSource_valid & _T_234; 
  assign cams_2_io_free_bits = io_d_tlSource_bits[2:0]; 
  assign cams_3_clock = clock; 
  assign cams_3_reset = reset; 
  assign cams_3_io_alloc_valid = _T_213 & extract_io_i_ready; 
  assign cams_3_io_alloc_bits = _T_6 ? _T_5 : _T_18; 
  assign cams_3_io_free_valid = io_d_tlSource_valid & _T_235; 
  assign cams_3_io_free_bits = io_d_tlSource_bits[2:0]; 
  assign cams_4_clock = clock; 
  assign cams_4_reset = reset; 
  assign cams_4_io_alloc_valid = _T_217 & extract_io_i_ready; 
  assign cams_4_io_alloc_bits = _T_6 ? _T_5 : _T_18; 
  assign cams_4_io_free_valid = io_d_tlSource_valid & _T_236; 
  assign cams_4_io_free_bits = io_d_tlSource_bits[2:0]; 
  assign cams_5_clock = clock; 
  assign cams_5_reset = reset; 
  assign cams_5_io_alloc_valid = _T_221 & extract_io_i_ready; 
  assign cams_5_io_alloc_bits = _T_6 ? _T_5 : _T_18; 
  assign cams_5_io_free_valid = io_d_tlSource_valid & _T_237; 
  assign cams_5_io_free_bits = io_d_tlSource_bits[2:0]; 
  assign cams_6_clock = clock; 
  assign cams_6_reset = reset; 
  assign cams_6_io_alloc_valid = _T_225 & extract_io_i_ready; 
  assign cams_6_io_alloc_bits = _T_6 ? _T_5 : _T_18; 
  assign cams_6_io_free_valid = io_d_tlSource_valid & _T_238; 
  assign cams_6_io_free_bits = io_d_tlSource_bits[2:0]; 
  assign cams_7_clock = clock; 
  assign cams_7_reset = reset; 
  assign cams_7_io_alloc_valid = _T_229 & extract_io_i_ready; 
  assign cams_7_io_alloc_bits = _T_6 ? _T_5 : _T_18; 
  assign cams_7_io_free_valid = io_d_tlSource_valid & _T_239; 
  assign cams_7_io_free_bits = io_d_tlSource_bits[2:0]; 
  assign extract_clock = clock; 
  assign extract_reset = reset; 
  assign extract_io_last = _T_72 | _T_74; 
  assign extract_io_i_valid = _T_185 & xmit; 
  assign extract_io_i_bits_opcode = _T_6 ? _T_1 : _T_10; 
  assign extract_io_i_bits_param = _T_6 ? _T_2 : _T_12; 
  assign extract_io_i_bits_size = _T_6 ? _T_3 : _T_14; 
  assign extract_io_i_bits_source = {_GEN_4,_GEN_23}; 
  assign extract_io_i_bits_address = _T_148[31:0]; 
  assign extract_io_i_bits_mask = {_T_180,_T_179}; 
  assign extract_io_i_bits_data = io_q_bits; 
  assign extract_io_o_ready = io_a_ready; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_10 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_12 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_14 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_16 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_18 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_20 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_22 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_23 = _RAND_8[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  a_first = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_143 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_75) begin
        if (_T_83) begin
          state <= 2'h1;
        end else begin
          if (_T_84) begin
            state <= 2'h2;
          end else begin
            if (_T_85) begin
              if (q_hasData) begin
                state <= 2'h3;
              end else begin
                state <= 2'h0;
              end
            end else begin
              if (_T_87) begin
                if (_T_88) begin
                  state <= 2'h3;
                end else begin
                  state <= 2'h0;
                end
              end
            end
          end
        end
      end
    end
    if (_T_6) begin
      _T_10 <= _T_1;
    end
    if (_T_6) begin
      _T_12 <= _T_2;
    end
    if (_T_6) begin
      _T_14 <= _T_3;
    end
    if (_T_6) begin
      _T_16 <= _T_4;
    end
    if (_T_6) begin
      _T_18 <= _T_5;
    end
    if (_T_19) begin
      _T_20 <= io_q_bits;
    end
    if (_T_21) begin
      _T_22 <= io_q_bits;
    end
    if (reset) begin
      _T_23 <= 11'h0;
    end else begin
      if (_T_75) begin
        if (_T_71) begin
          _T_23 <= _T_54;
        end else begin
          _T_23 <= _T_77;
        end
      end
    end
    if (_T_75) begin
      a_first <= _T_80;
    end
    if (a_first) begin
      if (3'h7 == _GEN_4) begin
        _T_143 <= _T_142_7;
      end else begin
        if (3'h6 == _GEN_4) begin
          _T_143 <= _T_142_6;
        end else begin
          if (3'h5 == _GEN_4) begin
            _T_143 <= _T_142_5;
          end else begin
            if (3'h4 == _GEN_4) begin
              _T_143 <= _T_142_4;
            end else begin
              if (3'h3 == _GEN_4) begin
                _T_143 <= _T_142_3;
              end else begin
                if (3'h2 == _GEN_4) begin
                  _T_143 <= _T_142_2;
                end else begin
                  if (3'h1 == _GEN_4) begin
                    _T_143 <= _T_142_1;
                  end else begin
                    _T_143 <= _T_142_0;
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module dual_SourceB( 
  input         clock, 
  input         reset, 
  output        io_bvalid, 
  output        io_q_ready, 
  input         io_q_valid, 
  input  [31:0] io_q_bits 
);
  wire  extract_clock; 
  wire  extract_reset; 
  wire  extract_io_last; 
  wire  extract_io_i_ready; 
  wire  extract_io_i_valid; 
  wire [2:0] extract_io_i_bits_opcode; 
  wire  extract_io_o_valid; 
  reg [1:0] state; 
  reg [31:0] _RAND_0;
  wire [2:0] _T_1; 
  wire [3:0] _T_3; 
  wire  _T_6; 
  reg [2:0] _T_10; 
  reg [31:0] _RAND_1;
  wire [2:0] _GEN_1; 
  reg [10:0] _T_25; 
  reg [31:0] _RAND_2;
  wire [15:0] _T_34; 
  wire [12:0] _T_35; 
  wire [9:0] _T_36; 
  wire  _T_37; 
  wire [10:0] _T_38; 
  wire [6:0] _T_43; 
  wire  _T_44; 
  wire [7:0] _T_45; 
  wire  _T_49; 
  wire  _T_50; 
  wire [10:0] _T_51; 
  wire [10:0] _T_53; 
  wire [7:0] _T_54; 
  wire [10:0] _GEN_15; 
  wire [10:0] _T_56; 
  wire  _T_73; 
  wire  _T_74; 
  wire  _T_75; 
  wire  _T_76; 
  wire  q_last; 
  wire  _T_77; 
  wire [10:0] _T_79; 
  wire  _T_81; 
  wire  q_hasData; 
  wire  _T_85; 
  wire  _T_86; 
  wire  _T_87; 
  wire  _T_89; 
  wire  _T_90; 
  wire  _T_126; 
  wire  xmit; 
  dual_ParitalExtractor_1 extract ( 
    .clock(extract_clock),
    .reset(extract_reset),
    .io_last(extract_io_last),
    .io_i_ready(extract_io_i_ready),
    .io_i_valid(extract_io_i_valid),
    .io_i_bits_opcode(extract_io_i_bits_opcode),
    .io_o_valid(extract_io_o_valid)
  );
  assign _T_1 = io_q_bits[5:3]; 
  assign _T_3 = io_q_bits[12:9]; 
  assign _T_6 = state == 2'h0; 
  assign _GEN_1 = _T_6 ? _T_1 : _T_10; 
  assign _T_34 = 16'h1 << _T_3; 
  assign _T_35 = _T_34[12:0]; 
  assign _T_36 = _T_35[12:3]; 
  assign _T_37 = _T_3 <= 4'h2; 
  assign _T_38 = {_T_36,_T_37}; 
  assign _T_43 = _T_35[12:6]; 
  assign _T_44 = _T_3 <= 4'h5; 
  assign _T_45 = {_T_43,_T_44}; 
  assign _T_49 = _T_1 == 3'h1; 
  assign _T_50 = _T_1[2]; 
  assign _T_51 = _T_50 ? 11'h0 : _T_38; 
  assign _T_53 = _T_51 + 11'h2; 
  assign _T_54 = _T_49 ? _T_45 : 8'h0; 
  assign _GEN_15 = {{3'd0}, _T_54}; 
  assign _T_56 = _T_53 + _GEN_15; 
  assign _T_73 = _T_25 == 11'h0; 
  assign _T_74 = _T_25 == 11'h1; 
  assign _T_75 = _T_56 == 11'h0; 
  assign _T_76 = _T_73 & _T_75; 
  assign q_last = _T_74 | _T_76; 
  assign _T_77 = io_q_ready & io_q_valid; 
  assign _T_79 = _T_25 - 11'h1; 
  assign _T_81 = _GEN_1[2]; 
  assign q_hasData = _T_81 == 1'h0; 
  assign _T_85 = 2'h0 == state; 
  assign _T_86 = 2'h1 == state; 
  assign _T_87 = 2'h2 == state; 
  assign _T_89 = 2'h3 == state; 
  assign _T_90 = q_last == 1'h0; 
  assign _T_126 = state == 2'h3; 
  assign xmit = q_last | _T_126; 
  assign io_bvalid = extract_io_o_valid; 
  assign io_q_ready = 1'h1; 
  assign extract_clock = clock; 
  assign extract_reset = reset; 
  assign extract_io_last = _T_74 | _T_76; 
  assign extract_io_i_valid = io_q_valid & xmit; 
  assign extract_io_i_bits_opcode = _T_6 ? _T_1 : _T_10; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_10 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[10:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_77) begin
        if (_T_85) begin
          state <= 2'h1;
        end else begin
          if (_T_86) begin
            state <= 2'h2;
          end else begin
            if (_T_87) begin
              if (q_hasData) begin
                state <= 2'h3;
              end else begin
                state <= 2'h0;
              end
            end else begin
              if (_T_89) begin
                if (_T_90) begin
                  state <= 2'h3;
                end else begin
                  state <= 2'h0;
                end
              end
            end
          end
        end
      end
    end
    if (_T_6) begin
      _T_10 <= _T_1;
    end
    if (reset) begin
      _T_25 <= 11'h0;
    end else begin
      if (_T_77) begin
        if (_T_73) begin
          _T_25 <= _T_56;
        end else begin
          _T_25 <= _T_79;
        end
      end
    end
  end
endmodule
module dual_SourceC( 
  input         clock, 
  input         reset, 
  input         io_c_ready, 
  output        io_c_valid, 
  output [2:0]  io_c_bits_opcode, 
  output [2:0]  io_c_bits_param, 
  output [3:0]  io_c_bits_size, 
  output [5:0]  io_c_bits_source, 
  output [31:0] io_c_bits_address, 
  output        io_q_ready, 
  input         io_q_valid, 
  input  [31:0] io_q_bits, 
  input         io_d_tlSource_valid, 
  input  [5:0]  io_d_tlSource_bits, 
  output [15:0] io_d_clSource 
);
  wire  cam_clock; 
  wire  cam_reset; 
  wire  cam_io_alloc_ready; 
  wire  cam_io_alloc_valid; 
  wire [15:0] cam_io_alloc_bits; 
  wire [2:0] cam_io_key; 
  wire  cam_io_free_valid; 
  wire [2:0] cam_io_free_bits; 
  wire [15:0] cam_io_data; 
  reg [1:0] state; 
  reg [31:0] _RAND_0;
  wire [2:0] _T_1; 
  wire [2:0] _T_2; 
  wire [3:0] _T_3; 
  wire [15:0] _T_5; 
  wire  _T_6; 
  reg [2:0] _T_10; 
  reg [31:0] _RAND_1;
  wire [2:0] _GEN_1; 
  reg [2:0] _T_12; 
  reg [31:0] _RAND_2;
  reg [3:0] _T_14; 
  reg [31:0] _RAND_3;
  reg [15:0] _T_19; 
  reg [31:0] _RAND_4;
  wire  _T_20; 
  reg [31:0] _T_21; 
  reg [31:0] _RAND_5;
  wire [31:0] _GEN_6; 
  wire  _T_22; 
  reg [31:0] _T_23; 
  reg [31:0] _RAND_6;
  wire [31:0] _GEN_7; 
  reg [10:0] _T_24; 
  reg [31:0] _RAND_7;
  wire [15:0] _T_33; 
  wire [12:0] _T_34; 
  wire [9:0] _T_35; 
  wire  _T_36; 
  wire [10:0] _T_37; 
  wire  _T_63; 
  wire [10:0] _T_64; 
  wire [10:0] _T_66; 
  wire  _T_72; 
  wire  _T_73; 
  wire  _T_74; 
  wire  _T_75; 
  wire  q_last; 
  wire  _T_76; 
  wire [10:0] _T_78; 
  wire  q_hasData; 
  wire  _T_80; 
  reg  c_first; 
  reg [31:0] _RAND_8;
  wire  _T_83; 
  wire  _T_84; 
  wire  _T_85; 
  wire  _T_87; 
  wire  _T_88; 
  wire [63:0] q_address; 
  wire [63:0] _T_90; 
  wire [64:0] _T_91; 
  wire [64:0] _T_92; 
  wire [64:0] _T_93; 
  wire  _T_94; 
  wire [63:0] _T_95; 
  wire [64:0] _T_96; 
  wire [64:0] _T_97; 
  wire [64:0] _T_98; 
  wire  _T_99; 
  wire [63:0] _T_100; 
  wire [64:0] _T_101; 
  wire [64:0] _T_102; 
  wire [64:0] _T_103; 
  wire  _T_104; 
  wire  _T_106; 
  wire  exists; 
  wire [64:0] _T_108; 
  wire [64:0] _T_125; 
  wire [64:0] _T_126; 
  wire  acquireOk; 
  wire  q_legal; 
  wire  _T_134; 
  wire  _T_135; 
  wire  q_release; 
  wire  _T_136; 
  wire  source_ok; 
  reg [2:0] _T_137; 
  reg [31:0] _RAND_9;
  wire [2:0] _GEN_15; 
  wire [2:0] _T_138; 
  wire [63:0] _T_139; 
  wire [35:0] _T_140; 
  wire [27:0] _T_141; 
  wire [63:0] _T_142; 
  wire  _T_143; 
  wire  stall; 
  wire  _T_144; 
  wire  xmit; 
  wire  _T_145; 
  wire  _T_146; 
  wire  _T_149; 
  wire  _T_150; 
  wire  _T_152; 
  wire  _T_153; 
  wire  _T_154; 
  dual_CAM cam ( 
    .clock(cam_clock),
    .reset(cam_reset),
    .io_alloc_ready(cam_io_alloc_ready),
    .io_alloc_valid(cam_io_alloc_valid),
    .io_alloc_bits(cam_io_alloc_bits),
    .io_key(cam_io_key),
    .io_free_valid(cam_io_free_valid),
    .io_free_bits(cam_io_free_bits),
    .io_data(cam_io_data)
  );
  assign _T_1 = io_q_bits[5:3]; 
  assign _T_2 = io_q_bits[8:6]; 
  assign _T_3 = io_q_bits[12:9]; 
  assign _T_5 = io_q_bits[31:16]; 
  assign _T_6 = state == 2'h0; 
  assign _GEN_1 = _T_6 ? _T_1 : _T_10; 
  assign _T_20 = state == 2'h1; 
  assign _GEN_6 = _T_20 ? io_q_bits : _T_21; 
  assign _T_22 = state == 2'h2; 
  assign _GEN_7 = _T_22 ? io_q_bits : _T_23; 
  assign _T_33 = 16'h1 << _T_3; 
  assign _T_34 = _T_33[12:0]; 
  assign _T_35 = _T_34[12:3]; 
  assign _T_36 = _T_3 <= 4'h2; 
  assign _T_37 = {_T_35,_T_36}; 
  assign _T_63 = _T_1[0]; 
  assign _T_64 = _T_63 ? _T_37 : 11'h0; 
  assign _T_66 = _T_64 + 11'h2; 
  assign _T_72 = _T_24 == 11'h0; 
  assign _T_73 = _T_24 == 11'h1; 
  assign _T_74 = _T_66 == 11'h0; 
  assign _T_75 = _T_72 & _T_74; 
  assign q_last = _T_73 | _T_75; 
  assign _T_76 = io_q_ready & io_q_valid; 
  assign _T_78 = _T_24 - 11'h1; 
  assign q_hasData = _GEN_1[0]; 
  assign _T_80 = state != 2'h3; 
  assign _T_83 = 2'h0 == state; 
  assign _T_84 = 2'h1 == state; 
  assign _T_85 = 2'h2 == state; 
  assign _T_87 = 2'h3 == state; 
  assign _T_88 = q_last == 1'h0; 
  assign q_address = {_GEN_7,_GEN_6}; 
  assign _T_90 = q_address ^ 64'h80000000; 
  assign _T_91 = {1'b0,$signed(_T_90)}; 
  assign _T_92 = $signed(_T_91) & $signed(-65'sh80000000); 
  assign _T_93 = $signed(_T_92); 
  assign _T_94 = $signed(_T_93) == $signed(65'sh0); 
  assign _T_95 = q_address ^ 64'h40000000; 
  assign _T_96 = {1'b0,$signed(_T_95)}; 
  assign _T_97 = $signed(_T_96) & $signed(-65'sh20000000); 
  assign _T_98 = $signed(_T_97); 
  assign _T_99 = $signed(_T_98) == $signed(65'sh0); 
  assign _T_100 = q_address ^ 64'h10000000; 
  assign _T_101 = {1'b0,$signed(_T_100)}; 
  assign _T_102 = $signed(_T_101) & $signed(-65'sh10000000); 
  assign _T_103 = $signed(_T_102); 
  assign _T_104 = $signed(_T_103) == $signed(65'sh0); 
  assign _T_106 = _T_94 | _T_99; 
  assign exists = _T_106 | _T_104; 
  assign _T_108 = {1'b0,$signed(q_address)}; 
  assign _T_125 = $signed(_T_108) & $signed(65'shc0000000); 
  assign _T_126 = $signed(_T_125); 
  assign acquireOk = $signed(_T_126) == $signed(65'sh0); 
  assign q_legal = exists & acquireOk; 
  assign _T_134 = _GEN_1 == 3'h6; 
  assign _T_135 = _GEN_1 == 3'h7; 
  assign q_release = _T_134 | _T_135; 
  assign _T_136 = q_release == 1'h0; 
  assign source_ok = _T_136 | cam_io_alloc_ready; 
  assign _GEN_15 = c_first ? cam_io_key : _T_137; 
  assign _T_138 = q_release ? _GEN_15 : 3'h0; 
  assign _T_139 = q_legal ? q_address : 64'h10000000; 
  assign _T_140 = _T_139[63:28]; 
  assign _T_141 = q_address[27:0]; 
  assign _T_142 = {_T_140,_T_141}; 
  assign _T_143 = source_ok == 1'h0; 
  assign stall = c_first & _T_143; 
  assign _T_144 = state == 2'h3; 
  assign xmit = q_last | _T_144; 
  assign _T_145 = stall == 1'h0; 
  assign _T_146 = io_q_valid & _T_145; 
  assign _T_149 = io_c_ready & _T_145; 
  assign _T_150 = xmit == 1'h0; 
  assign _T_152 = q_release & c_first; 
  assign _T_153 = _T_152 & xmit; 
  assign _T_154 = _T_153 & io_q_valid; 
  assign io_c_valid = _T_146 & xmit; 
  assign io_c_bits_opcode = _T_6 ? _T_1 : _T_10; 
  assign io_c_bits_param = _T_6 ? _T_2 : _T_12; 
  assign io_c_bits_size = _T_6 ? _T_3 : _T_14; 
  assign io_c_bits_source = {{3'd0}, _T_138}; 
  assign io_c_bits_address = _T_142[31:0]; 
  assign io_q_ready = _T_149 | _T_150; 
  assign io_d_clSource = cam_io_data; 
  assign cam_clock = clock; 
  assign cam_reset = reset; 
  assign cam_io_alloc_valid = _T_154 & io_c_ready; 
  assign cam_io_alloc_bits = _T_6 ? _T_5 : _T_19; 
  assign cam_io_free_valid = io_d_tlSource_valid; 
  assign cam_io_free_bits = io_d_tlSource_bits[2:0]; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_10 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_12 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_14 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_19 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_21 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_23 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_24 = _RAND_7[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  c_first = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_137 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_76) begin
        if (_T_83) begin
          state <= 2'h1;
        end else begin
          if (_T_84) begin
            state <= 2'h2;
          end else begin
            if (_T_85) begin
              if (q_hasData) begin
                state <= 2'h3;
              end else begin
                state <= 2'h0;
              end
            end else begin
              if (_T_87) begin
                if (_T_88) begin
                  state <= 2'h3;
                end else begin
                  state <= 2'h0;
                end
              end
            end
          end
        end
      end
    end
    if (_T_6) begin
      _T_10 <= _T_1;
    end
    if (_T_6) begin
      _T_12 <= _T_2;
    end
    if (_T_6) begin
      _T_14 <= _T_3;
    end
    if (_T_6) begin
      _T_19 <= _T_5;
    end
    if (_T_20) begin
      _T_21 <= io_q_bits;
    end
    if (_T_22) begin
      _T_23 <= io_q_bits;
    end
    if (reset) begin
      _T_24 <= 11'h0;
    end else begin
      if (_T_76) begin
        if (_T_72) begin
          _T_24 <= _T_66;
        end else begin
          _T_24 <= _T_78;
        end
      end
    end
    if (_T_76) begin
      c_first <= _T_80;
    end
    if (c_first) begin
      _T_137 <= cam_io_key;
    end
  end
endmodule
module dual_SourceD( 
  input         clock, 
  input         reset, 
  input         io_d_ready, 
  output        io_d_valid, 
  output [2:0]  io_d_bits_opcode, 
  output [1:0]  io_d_bits_param, 
  output [2:0]  io_d_bits_size, 
  output [2:0]  io_d_bits_source, 
  output [4:0]  io_d_bits_sink, 
  output        io_d_bits_denied, 
  output [31:0] io_d_bits_data, 
  output        io_d_bits_corrupt, 
  output        io_q_ready, 
  input         io_q_valid, 
  input  [31:0] io_q_bits, 
  output [15:0] io_e_clSink 
);
  wire  cam_clock; 
  wire  cam_reset; 
  wire  cam_io_alloc_ready; 
  wire  cam_io_alloc_valid; 
  wire [15:0] cam_io_alloc_bits; 
  wire [4:0] cam_io_key; 
  wire [15:0] cam_io_data; 
  reg [1:0] state; 
  reg [31:0] _RAND_0;
  wire [2:0] _T_1; 
  wire [2:0] _T_2; 
  wire [3:0] _T_3; 
  wire [2:0] _T_4; 
  wire [15:0] _T_5; 
  wire  _T_6; 
  reg [2:0] _T_10; 
  reg [31:0] _RAND_1;
  wire [2:0] _GEN_1; 
  reg [2:0] _T_12; 
  reg [31:0] _RAND_2;
  wire [2:0] _GEN_2; 
  reg [3:0] _T_14; 
  reg [31:0] _RAND_3;
  wire [3:0] _GEN_3; 
  reg [2:0] _T_16; 
  reg [31:0] _RAND_4;
  wire [2:0] _GEN_4; 
  reg [15:0] _T_18; 
  reg [31:0] _RAND_5;
  wire [15:0] _GEN_5; 
  wire [15:0] _T_19; 
  wire  _T_20; 
  reg [15:0] _T_21; 
  reg [31:0] _RAND_6;
  wire  _T_22; 
  wire  _T_23; 
  wire  q_grant; 
  reg [10:0] _T_24; 
  reg [31:0] _RAND_7;
  wire [15:0] _T_33; 
  wire [12:0] _T_34; 
  wire [9:0] _T_35; 
  wire  _T_36; 
  wire [10:0] _T_37; 
  wire  _T_45; 
  wire  _T_46; 
  wire  _T_47; 
  wire  _T_63; 
  wire [10:0] _T_64; 
  wire [10:0] _GEN_32; 
  wire [10:0] _T_70; 
  wire  _T_72; 
  wire  _T_73; 
  wire  _T_74; 
  wire  _T_75; 
  wire  q_last; 
  wire  _T_76; 
  wire [10:0] _T_78; 
  wire  _T_80; 
  reg  d_first; 
  reg [31:0] _RAND_8;
  wire  _T_83; 
  wire  _T_85; 
  wire  _T_86; 
  wire  _T_87; 
  wire  sink_ok; 
  reg [4:0] _T_88; 
  reg [31:0] _RAND_9;
  wire [4:0] _GEN_13; 
  wire  _T_89; 
  wire  stall; 
  wire  _T_90; 
  wire  xmit; 
  wire [1:0] _T_92; 
  wire [1:0] _GEN_15; 
  wire [1:0] _GEN_16; 
  wire [1:0] _GEN_17; 
  wire [2:0] _GEN_19; 
  wire [2:0] _GEN_20; 
  wire [2:0] _GEN_21; 
  wire [2:0] _T_94_1; 
  wire [2:0] _GEN_23; 
  wire [2:0] _GEN_24; 
  wire [2:0] _GEN_25; 
  wire [2:0] _GEN_26; 
  wire [2:0] _GEN_27; 
  wire [2:0] _GEN_28; 
  wire  _T_97; 
  wire  _T_99; 
  wire  _T_100; 
  wire  _T_103; 
  wire  _T_104; 
  wire  _T_106; 
  wire  _T_107; 
  wire  _T_108; 
  dual_CAM_9 cam ( 
    .clock(cam_clock),
    .reset(cam_reset),
    .io_alloc_ready(cam_io_alloc_ready),
    .io_alloc_valid(cam_io_alloc_valid),
    .io_alloc_bits(cam_io_alloc_bits),
    .io_key(cam_io_key),
    .io_data(cam_io_data)
  );
  assign _T_1 = io_q_bits[5:3]; 
  assign _T_2 = io_q_bits[8:6]; 
  assign _T_3 = io_q_bits[12:9]; 
  assign _T_4 = io_q_bits[15:13]; 
  assign _T_5 = io_q_bits[31:16]; 
  assign _T_6 = state == 2'h0; 
  assign _GEN_1 = _T_6 ? _T_1 : _T_10; 
  assign _GEN_2 = _T_6 ? _T_2 : _T_12; 
  assign _GEN_3 = _T_6 ? _T_3 : _T_14; 
  assign _GEN_4 = _T_6 ? _T_4 : _T_16; 
  assign _GEN_5 = _T_6 ? _T_5 : _T_18; 
  assign _T_19 = io_q_bits[15:0]; 
  assign _T_20 = state == 2'h1; 
  assign _T_22 = _GEN_1 == 3'h4; 
  assign _T_23 = _GEN_1 == 3'h5; 
  assign q_grant = _T_22 | _T_23; 
  assign _T_33 = 16'h1 << _T_3; 
  assign _T_34 = _T_33[12:0]; 
  assign _T_35 = _T_34[12:3]; 
  assign _T_36 = _T_3 <= 4'h2; 
  assign _T_37 = {_T_35,_T_36}; 
  assign _T_45 = _T_1 == 3'h4; 
  assign _T_46 = _T_1 == 3'h5; 
  assign _T_47 = _T_45 | _T_46; 
  assign _T_63 = _T_1[0]; 
  assign _T_64 = _T_63 ? _T_37 : 11'h0; 
  assign _GEN_32 = {{10'd0}, _T_47}; 
  assign _T_70 = _T_64 + _GEN_32; 
  assign _T_72 = _T_24 == 11'h0; 
  assign _T_73 = _T_24 == 11'h1; 
  assign _T_74 = _T_70 == 11'h0; 
  assign _T_75 = _T_72 & _T_74; 
  assign q_last = _T_73 | _T_75; 
  assign _T_76 = io_q_ready & io_q_valid; 
  assign _T_78 = _T_24 - 11'h1; 
  assign _T_80 = state != 2'h2; 
  assign _T_83 = 2'h0 == state; 
  assign _T_85 = 2'h1 == state; 
  assign _T_86 = 2'h2 == state; 
  assign _T_87 = q_grant == 1'h0; 
  assign sink_ok = _T_87 | cam_io_alloc_ready; 
  assign _GEN_13 = d_first ? cam_io_key : _T_88; 
  assign _T_89 = sink_ok == 1'h0; 
  assign stall = d_first & _T_89; 
  assign _T_90 = state == 2'h2; 
  assign xmit = q_last | _T_90; 
  assign _T_92 = _GEN_5[1:0]; 
  assign _GEN_15 = 2'h1 == _T_92 ? 2'h1 : 2'h0; 
  assign _GEN_16 = 2'h2 == _T_92 ? 2'h2 : _GEN_15; 
  assign _GEN_17 = 2'h3 == _T_92 ? 2'h3 : _GEN_16; 
  assign _GEN_19 = 2'h1 == _T_92 ? 3'h5 : 3'h4; 
  assign _GEN_20 = 2'h2 == _T_92 ? 3'h6 : _GEN_19; 
  assign _GEN_21 = 2'h3 == _T_92 ? 3'h7 : _GEN_20; 
  assign _T_94_1 = {{1'd0}, _GEN_17}; 
  assign _GEN_23 = 3'h1 == _GEN_4 ? _T_94_1 : 3'h0; 
  assign _GEN_24 = 3'h2 == _GEN_4 ? _GEN_21 : _GEN_23; 
  assign _GEN_25 = 3'h3 == _GEN_4 ? 3'h0 : _GEN_24; 
  assign _GEN_26 = 3'h4 == _GEN_4 ? 3'h0 : _GEN_25; 
  assign _GEN_27 = 3'h5 == _GEN_4 ? 3'h0 : _GEN_26; 
  assign _GEN_28 = 3'h6 == _GEN_4 ? 3'h0 : _GEN_27; 
  assign _T_97 = io_d_bits_opcode[0]; 
  assign _T_99 = stall == 1'h0; 
  assign _T_100 = io_q_valid & _T_99; 
  assign _T_103 = io_d_ready & _T_99; 
  assign _T_104 = xmit == 1'h0; 
  assign _T_106 = q_grant & d_first; 
  assign _T_107 = _T_106 & xmit; 
  assign _T_108 = _T_107 & io_q_valid; 
  assign io_d_valid = _T_100 & xmit; 
  assign io_d_bits_opcode = _T_6 ? _T_1 : _T_10; 
  assign io_d_bits_param = _GEN_2[1:0]; 
  assign io_d_bits_size = _GEN_3[2:0]; 
  assign io_d_bits_source = 3'h7 == _GEN_4 ? 3'h0 : _GEN_28; 
  assign io_d_bits_sink = q_grant ? _GEN_13 : 5'h0; 
  assign io_d_bits_denied = _GEN_2[2:2]; 
  assign io_d_bits_data = io_q_bits; 
  assign io_d_bits_corrupt = io_d_bits_denied & _T_97; 
  assign io_q_ready = _T_103 | _T_104; 
  assign io_e_clSink = cam_io_data; 
  assign cam_clock = clock; 
  assign cam_reset = reset; 
  assign cam_io_alloc_valid = _T_108 & io_d_ready; 
  assign cam_io_alloc_bits = _T_20 ? _T_19 : _T_21; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_10 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_12 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_14 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_16 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_18 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_21 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_24 = _RAND_7[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  d_first = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_88 = _RAND_9[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_76) begin
        if (_T_83) begin
          if (q_grant) begin
            state <= 2'h1;
          end else begin
            if (q_last) begin
              state <= 2'h0;
            end else begin
              state <= 2'h2;
            end
          end
        end else begin
          if (_T_85) begin
            if (q_last) begin
              state <= 2'h0;
            end else begin
              state <= 2'h2;
            end
          end else begin
            if (_T_86) begin
              if (q_last) begin
                state <= 2'h0;
              end else begin
                state <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (_T_6) begin
      _T_10 <= _T_1;
    end
    if (_T_6) begin
      _T_12 <= _T_2;
    end
    if (_T_6) begin
      _T_14 <= _T_3;
    end
    if (_T_6) begin
      _T_16 <= _T_4;
    end
    if (_T_6) begin
      _T_18 <= _T_5;
    end
    if (_T_20) begin
      _T_21 <= _T_19;
    end
    if (reset) begin
      _T_24 <= 11'h0;
    end else begin
      if (_T_76) begin
        if (_T_72) begin
          _T_24 <= _T_70;
        end else begin
          _T_24 <= _T_78;
        end
      end
    end
    if (_T_76) begin
      d_first <= _T_80;
    end
    if (d_first) begin
      _T_88 <= cam_io_key;
    end
  end
endmodule
module dual_SourceE( 
  input         io_e_ready, 
  output        io_e_valid, 
  output        io_e_bits_sink, 
  output        io_q_ready, 
  input         io_q_valid, 
  input  [31:0] io_q_bits 
);
  wire [15:0] q_sink; 
  assign q_sink = io_q_bits[31:16]; 
  assign io_e_valid = io_q_valid; 
  assign io_e_bits_sink = q_sink[0]; 
  assign io_q_ready = io_e_ready; 
endmodule
module dual_SynchronizerShiftReg_w100_d1( 
  input         clock, 
  input  [99:0] io_d, 
  output [99:0] io_q 
);
  reg [99:0] sync_0; 
  reg [127:0] _RAND_0;
  assign io_q = sync_0; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  sync_0 = _RAND_0[99:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    sync_0 <= io_d;
  end
endmodule
module dual_SynchronizerShiftReg_w32_d1( 
  input         clock, 
  input  [31:0] io_d, 
  output [31:0] io_q 
);
  reg [31:0] sync_0; 
  reg [31:0] _RAND_0;
  assign io_q = sync_0; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sync_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    sync_0 <= io_d;
  end
endmodule
module dual_TLAtomicAutomata( 
  input         clock, 
  input         reset, 
  output        auto_in_a_ready, 
  input         auto_in_a_valid, 
  input  [2:0]  auto_in_a_bits_opcode, 
  input  [2:0]  auto_in_a_bits_param, 
  input  [3:0]  auto_in_a_bits_size, 
  input  [6:0]  auto_in_a_bits_source, 
  input  [31:0] auto_in_a_bits_address, 
  input  [7:0]  auto_in_a_bits_mask, 
  input  [63:0] auto_in_a_bits_data, 
  output        auto_in_c_ready, 
  input         auto_in_c_valid, 
  input  [2:0]  auto_in_c_bits_opcode, 
  input  [2:0]  auto_in_c_bits_param, 
  input  [3:0]  auto_in_c_bits_size, 
  input  [6:0]  auto_in_c_bits_source, 
  input  [31:0] auto_in_c_bits_address, 
  input         auto_in_c_bits_corrupt, 
  input         auto_in_d_ready, 
  output        auto_in_d_valid, 
  output [2:0]  auto_in_d_bits_opcode, 
  output [1:0]  auto_in_d_bits_param, 
  output [3:0]  auto_in_d_bits_size, 
  output [6:0]  auto_in_d_bits_source, 
  output        auto_in_d_bits_sink, 
  output        auto_in_d_bits_denied, 
  output [63:0] auto_in_d_bits_data, 
  output        auto_in_d_bits_corrupt, 
  output        auto_in_e_ready, 
  input         auto_in_e_valid, 
  input         auto_in_e_bits_sink, 
  input         auto_out_a_ready, 
  output        auto_out_a_valid, 
  output [2:0]  auto_out_a_bits_opcode, 
  output [2:0]  auto_out_a_bits_param, 
  output [3:0]  auto_out_a_bits_size, 
  output [6:0]  auto_out_a_bits_source, 
  output [31:0] auto_out_a_bits_address, 
  output [7:0]  auto_out_a_bits_mask, 
  output [63:0] auto_out_a_bits_data, 
  output        auto_out_a_bits_corrupt, 
  input         auto_out_c_ready, 
  output        auto_out_c_valid, 
  output [2:0]  auto_out_c_bits_opcode, 
  output [2:0]  auto_out_c_bits_param, 
  output [3:0]  auto_out_c_bits_size, 
  output [6:0]  auto_out_c_bits_source, 
  output [31:0] auto_out_c_bits_address, 
  output        auto_out_c_bits_corrupt, 
  output        auto_out_d_ready, 
  input         auto_out_d_valid, 
  input  [2:0]  auto_out_d_bits_opcode, 
  input  [1:0]  auto_out_d_bits_param, 
  input  [3:0]  auto_out_d_bits_size, 
  input  [6:0]  auto_out_d_bits_source, 
  input         auto_out_d_bits_sink, 
  input         auto_out_d_bits_denied, 
  input  [63:0] auto_out_d_bits_data, 
  input         auto_out_d_bits_corrupt, 
  input         auto_out_e_ready, 
  output        auto_out_e_valid, 
  output        auto_out_e_bits_sink 
);
  wire  TLMonitor_clock; 
  wire  TLMonitor_reset; 
  wire  TLMonitor_io_in_a_ready; 
  wire  TLMonitor_io_in_a_valid; 
  wire [2:0] TLMonitor_io_in_a_bits_opcode; 
  wire [2:0] TLMonitor_io_in_a_bits_param; 
  wire [3:0] TLMonitor_io_in_a_bits_size; 
  wire [6:0] TLMonitor_io_in_a_bits_source; 
  wire [31:0] TLMonitor_io_in_a_bits_address; 
  wire [7:0] TLMonitor_io_in_a_bits_mask; 
  wire  TLMonitor_io_in_c_ready; 
  wire  TLMonitor_io_in_c_valid; 
  wire [2:0] TLMonitor_io_in_c_bits_opcode; 
  wire [2:0] TLMonitor_io_in_c_bits_param; 
  wire [3:0] TLMonitor_io_in_c_bits_size; 
  wire [6:0] TLMonitor_io_in_c_bits_source; 
  wire [31:0] TLMonitor_io_in_c_bits_address; 
  wire  TLMonitor_io_in_c_bits_corrupt; 
  wire  TLMonitor_io_in_d_ready; 
  wire  TLMonitor_io_in_d_valid; 
  wire [2:0] TLMonitor_io_in_d_bits_opcode; 
  wire [1:0] TLMonitor_io_in_d_bits_param; 
  wire [3:0] TLMonitor_io_in_d_bits_size; 
  wire [6:0] TLMonitor_io_in_d_bits_source; 
  wire  TLMonitor_io_in_d_bits_sink; 
  wire  TLMonitor_io_in_d_bits_denied; 
  wire  TLMonitor_io_in_d_bits_corrupt; 
  wire  TLMonitor_io_in_e_ready; 
  wire  TLMonitor_io_in_e_valid; 
  wire  TLMonitor_io_in_e_bits_sink; 
  reg [1:0] _T_10_0_state; 
  reg [31:0] _RAND_0;
  reg [2:0] _T_11_0_bits_opcode; 
  reg [31:0] _RAND_1;
  reg [2:0] _T_11_0_bits_param; 
  reg [31:0] _RAND_2;
  reg [3:0] _T_11_0_bits_size; 
  reg [31:0] _RAND_3;
  reg [6:0] _T_11_0_bits_source; 
  reg [31:0] _RAND_4;
  reg [31:0] _T_11_0_bits_address; 
  reg [31:0] _RAND_5;
  reg [7:0] _T_11_0_bits_mask; 
  reg [31:0] _RAND_6;
  reg [63:0] _T_11_0_bits_data; 
  reg [63:0] _RAND_7;
  reg [1:0] _T_11_0_fifoId; 
  reg [31:0] _RAND_8;
  reg [3:0] _T_11_0_lut; 
  reg [31:0] _RAND_9;
  reg [63:0] _T_12_0_data; 
  reg [63:0] _RAND_10;
  reg  _T_12_0_denied; 
  reg [31:0] _RAND_11;
  reg  _T_12_0_corrupt; 
  reg [31:0] _RAND_12;
  wire  _T_13; 
  wire  _T_14; 
  wire  _T_15; 
  wire  _T_17; 
  wire  _T_18; 
  wire [31:0] _T_25; 
  wire [32:0] _T_26; 
  wire [32:0] _T_27; 
  wire [32:0] _T_28; 
  wire  _T_29; 
  wire [32:0] _T_37; 
  wire [32:0] _T_38; 
  wire [32:0] _T_39; 
  wire  _T_40; 
  wire  _T_71; 
  wire  _T_72; 
  wire  _T_73; 
  wire  _T_74; 
  wire [1:0] _T_95; 
  wire [1:0] _GEN_43; 
  wire [1:0] _T_97; 
  wire  _T_99; 
  wire  _T_100; 
  wire  _T_104; 
  wire  _T_105; 
  wire [1:0] _T_106; 
  wire  _T_107; 
  wire  _T_108; 
  wire [1:0] _T_109; 
  wire  _T_110; 
  wire  _T_111; 
  wire [1:0] _T_112; 
  wire  _T_113; 
  wire  _T_114; 
  wire [1:0] _T_115; 
  wire  _T_116; 
  wire  _T_117; 
  wire [1:0] _T_118; 
  wire  _T_119; 
  wire  _T_120; 
  wire [1:0] _T_121; 
  wire  _T_122; 
  wire  _T_123; 
  wire [1:0] _T_124; 
  wire  _T_125; 
  wire  _T_126; 
  wire [1:0] _T_127; 
  wire  _T_128; 
  wire  _T_129; 
  wire [1:0] _T_130; 
  wire  _T_131; 
  wire  _T_132; 
  wire [1:0] _T_133; 
  wire  _T_134; 
  wire  _T_135; 
  wire [1:0] _T_136; 
  wire  _T_137; 
  wire  _T_138; 
  wire [1:0] _T_139; 
  wire  _T_140; 
  wire  _T_141; 
  wire [1:0] _T_142; 
  wire  _T_143; 
  wire  _T_144; 
  wire [1:0] _T_145; 
  wire  _T_146; 
  wire  _T_147; 
  wire [1:0] _T_148; 
  wire  _T_149; 
  wire  _T_150; 
  wire [1:0] _T_151; 
  wire  _T_152; 
  wire  _T_153; 
  wire [1:0] _T_154; 
  wire  _T_155; 
  wire  _T_156; 
  wire [1:0] _T_157; 
  wire  _T_158; 
  wire  _T_159; 
  wire [1:0] _T_160; 
  wire  _T_161; 
  wire  _T_162; 
  wire [1:0] _T_163; 
  wire  _T_164; 
  wire  _T_165; 
  wire [1:0] _T_166; 
  wire  _T_167; 
  wire  _T_168; 
  wire [1:0] _T_169; 
  wire  _T_170; 
  wire  _T_171; 
  wire [1:0] _T_172; 
  wire  _T_173; 
  wire  _T_174; 
  wire [1:0] _T_175; 
  wire  _T_176; 
  wire  _T_177; 
  wire [1:0] _T_178; 
  wire  _T_179; 
  wire  _T_180; 
  wire [1:0] _T_181; 
  wire  _T_182; 
  wire  _T_183; 
  wire [1:0] _T_184; 
  wire  _T_185; 
  wire  _T_186; 
  wire [1:0] _T_187; 
  wire  _T_188; 
  wire  _T_189; 
  wire [1:0] _T_190; 
  wire  _T_191; 
  wire  _T_192; 
  wire [1:0] _T_193; 
  wire  _T_194; 
  wire  _T_195; 
  wire [1:0] _T_196; 
  wire  _T_197; 
  wire  _T_198; 
  wire [1:0] _T_199; 
  wire  _T_200; 
  wire  _T_201; 
  wire [1:0] _T_202; 
  wire  _T_203; 
  wire  _T_204; 
  wire [1:0] _T_205; 
  wire  _T_206; 
  wire  _T_207; 
  wire [1:0] _T_208; 
  wire  _T_209; 
  wire  _T_210; 
  wire [1:0] _T_211; 
  wire  _T_212; 
  wire  _T_213; 
  wire [1:0] _T_214; 
  wire  _T_215; 
  wire  _T_216; 
  wire [1:0] _T_217; 
  wire  _T_218; 
  wire  _T_219; 
  wire [1:0] _T_220; 
  wire  _T_221; 
  wire  _T_222; 
  wire [1:0] _T_223; 
  wire  _T_224; 
  wire  _T_225; 
  wire [1:0] _T_226; 
  wire  _T_227; 
  wire  _T_228; 
  wire [1:0] _T_229; 
  wire  _T_230; 
  wire  _T_231; 
  wire [1:0] _T_232; 
  wire  _T_233; 
  wire  _T_234; 
  wire [1:0] _T_235; 
  wire  _T_236; 
  wire  _T_237; 
  wire [1:0] _T_238; 
  wire  _T_239; 
  wire  _T_240; 
  wire [1:0] _T_241; 
  wire  _T_242; 
  wire  _T_243; 
  wire [1:0] _T_244; 
  wire  _T_245; 
  wire  _T_246; 
  wire [1:0] _T_247; 
  wire  _T_248; 
  wire  _T_249; 
  wire [1:0] _T_250; 
  wire  _T_251; 
  wire  _T_252; 
  wire [1:0] _T_253; 
  wire  _T_254; 
  wire  _T_255; 
  wire [1:0] _T_256; 
  wire  _T_257; 
  wire  _T_258; 
  wire [1:0] _T_259; 
  wire  _T_260; 
  wire  _T_261; 
  wire [1:0] _T_262; 
  wire  _T_263; 
  wire  _T_264; 
  wire [1:0] _T_265; 
  wire  _T_266; 
  wire  _T_267; 
  wire [1:0] _T_268; 
  wire  _T_269; 
  wire  _T_270; 
  wire [1:0] _T_271; 
  wire  _T_272; 
  wire  _T_273; 
  wire [1:0] _T_274; 
  wire  _T_275; 
  wire  _T_276; 
  wire [1:0] _T_277; 
  wire  _T_278; 
  wire  _T_279; 
  wire [1:0] _T_280; 
  wire  _T_281; 
  wire  _T_282; 
  wire [1:0] _T_283; 
  wire  _T_284; 
  wire  _T_285; 
  wire [1:0] _T_286; 
  wire  _T_287; 
  wire  _T_288; 
  wire [1:0] _T_289; 
  wire  _T_290; 
  wire  _T_291; 
  wire [1:0] _T_292; 
  wire  _T_293; 
  wire  _T_294; 
  wire [1:0] _T_295; 
  wire [3:0] _T_296; 
  wire  _T_297; 
  wire [3:0] _T_298; 
  wire  _T_299; 
  wire [3:0] _T_300; 
  wire  _T_301; 
  wire [3:0] _T_302; 
  wire  _T_303; 
  wire [3:0] _T_304; 
  wire  _T_305; 
  wire [3:0] _T_306; 
  wire  _T_307; 
  wire [3:0] _T_308; 
  wire  _T_309; 
  wire [3:0] _T_310; 
  wire  _T_311; 
  wire [3:0] _T_312; 
  wire  _T_313; 
  wire [3:0] _T_314; 
  wire  _T_315; 
  wire [3:0] _T_316; 
  wire  _T_317; 
  wire [3:0] _T_318; 
  wire  _T_319; 
  wire [3:0] _T_320; 
  wire  _T_321; 
  wire [3:0] _T_322; 
  wire  _T_323; 
  wire [3:0] _T_324; 
  wire  _T_325; 
  wire [3:0] _T_326; 
  wire  _T_327; 
  wire [3:0] _T_328; 
  wire  _T_329; 
  wire [3:0] _T_330; 
  wire  _T_331; 
  wire [3:0] _T_332; 
  wire  _T_333; 
  wire [3:0] _T_334; 
  wire  _T_335; 
  wire [3:0] _T_336; 
  wire  _T_337; 
  wire [3:0] _T_338; 
  wire  _T_339; 
  wire [3:0] _T_340; 
  wire  _T_341; 
  wire [3:0] _T_342; 
  wire  _T_343; 
  wire [3:0] _T_344; 
  wire  _T_345; 
  wire [3:0] _T_346; 
  wire  _T_347; 
  wire [3:0] _T_348; 
  wire  _T_349; 
  wire [3:0] _T_350; 
  wire  _T_351; 
  wire [3:0] _T_352; 
  wire  _T_353; 
  wire [3:0] _T_354; 
  wire  _T_355; 
  wire [3:0] _T_356; 
  wire  _T_357; 
  wire [3:0] _T_358; 
  wire  _T_359; 
  wire [3:0] _T_360; 
  wire  _T_361; 
  wire [3:0] _T_362; 
  wire  _T_363; 
  wire [3:0] _T_364; 
  wire  _T_365; 
  wire [3:0] _T_366; 
  wire  _T_367; 
  wire [3:0] _T_368; 
  wire  _T_369; 
  wire [3:0] _T_370; 
  wire  _T_371; 
  wire [3:0] _T_372; 
  wire  _T_373; 
  wire [3:0] _T_374; 
  wire  _T_375; 
  wire [3:0] _T_376; 
  wire  _T_377; 
  wire [3:0] _T_378; 
  wire  _T_379; 
  wire [3:0] _T_380; 
  wire  _T_381; 
  wire [3:0] _T_382; 
  wire  _T_383; 
  wire [3:0] _T_384; 
  wire  _T_385; 
  wire [3:0] _T_386; 
  wire  _T_387; 
  wire [3:0] _T_388; 
  wire  _T_389; 
  wire [3:0] _T_390; 
  wire  _T_391; 
  wire [3:0] _T_392; 
  wire  _T_393; 
  wire [3:0] _T_394; 
  wire  _T_395; 
  wire [3:0] _T_396; 
  wire  _T_397; 
  wire [3:0] _T_398; 
  wire  _T_399; 
  wire [3:0] _T_400; 
  wire  _T_401; 
  wire [3:0] _T_402; 
  wire  _T_403; 
  wire [3:0] _T_404; 
  wire  _T_405; 
  wire [3:0] _T_406; 
  wire  _T_407; 
  wire [3:0] _T_408; 
  wire  _T_409; 
  wire [3:0] _T_410; 
  wire  _T_411; 
  wire [3:0] _T_412; 
  wire  _T_413; 
  wire [3:0] _T_414; 
  wire  _T_415; 
  wire [3:0] _T_416; 
  wire  _T_417; 
  wire [3:0] _T_418; 
  wire  _T_419; 
  wire [3:0] _T_420; 
  wire  _T_421; 
  wire [3:0] _T_422; 
  wire  _T_423; 
  wire [7:0] _T_430; 
  wire [15:0] _T_438; 
  wire [7:0] _T_445; 
  wire [31:0] _T_454; 
  wire [7:0] _T_461; 
  wire [15:0] _T_469; 
  wire [7:0] _T_476; 
  wire [31:0] _T_485; 
  wire [63:0] _T_486; 
  wire  _T_487; 
  wire  _T_488; 
  wire  _T_489; 
  wire [7:0] _T_490; 
  wire [6:0] _T_491; 
  wire [7:0] _GEN_44; 
  wire [7:0] _T_492; 
  wire [7:0] _T_493; 
  wire [7:0] _T_508; 
  wire [7:0] _T_523; 
  wire [7:0] _T_524; 
  wire [8:0] _T_525; 
  wire [7:0] _T_526; 
  wire [7:0] _T_527; 
  wire [8:0] _T_528; 
  wire [7:0] _T_529; 
  wire [8:0] _T_530; 
  wire [7:0] _T_531; 
  wire [7:0] _T_532; 
  wire [9:0] _T_533; 
  wire [7:0] _T_534; 
  wire [7:0] _T_535; 
  wire [11:0] _T_536; 
  wire [7:0] _T_537; 
  wire [7:0] _T_538; 
  wire  _T_540; 
  wire  _T_541; 
  wire  _T_542; 
  wire  _T_543; 
  wire  _T_544; 
  wire  _T_545; 
  wire  _T_546; 
  wire  _T_547; 
  wire [7:0] _T_549; 
  wire [7:0] _T_551; 
  wire [7:0] _T_553; 
  wire [7:0] _T_555; 
  wire [7:0] _T_557; 
  wire [7:0] _T_559; 
  wire [7:0] _T_561; 
  wire [7:0] _T_563; 
  wire [63:0] _T_570; 
  wire [8:0] _T_571; 
  wire [7:0] _T_572; 
  wire [7:0] _T_573; 
  wire [9:0] _T_574; 
  wire [7:0] _T_575; 
  wire [7:0] _T_576; 
  wire [11:0] _T_577; 
  wire [7:0] _T_578; 
  wire [7:0] _T_579; 
  wire  _T_581; 
  wire  _T_582; 
  wire  _T_583; 
  wire  _T_584; 
  wire  _T_585; 
  wire  _T_586; 
  wire  _T_587; 
  wire  _T_588; 
  wire [7:0] _T_590; 
  wire [7:0] _T_592; 
  wire [7:0] _T_594; 
  wire [7:0] _T_596; 
  wire [7:0] _T_598; 
  wire [7:0] _T_600; 
  wire [7:0] _T_602; 
  wire [7:0] _T_604; 
  wire [63:0] _T_611; 
  wire  _T_612; 
  wire  _T_613; 
  wire  _T_614; 
  wire  _T_615; 
  wire  _T_616; 
  wire  _T_617; 
  wire  _T_618; 
  wire  _T_619; 
  wire [7:0] _T_621; 
  wire [7:0] _T_623; 
  wire [7:0] _T_625; 
  wire [7:0] _T_627; 
  wire [7:0] _T_629; 
  wire [7:0] _T_631; 
  wire [7:0] _T_633; 
  wire [7:0] _T_635; 
  wire [63:0] _T_642; 
  wire [63:0] _T_643; 
  wire [63:0] _T_644; 
  wire [63:0] _T_645; 
  wire [63:0] _T_646; 
  wire [63:0] _T_647; 
  wire [63:0] _T_648; 
  wire [63:0] _T_650; 
  wire  _T_651; 
  wire  _T_652; 
  wire  _T_654; 
  wire  _T_655; 
  wire  _T_656; 
  wire  _T_657; 
  wire  _T_658; 
  wire  _T_659; 
  wire [63:0] _T_660; 
  wire [63:0] _T_661; 
  wire  _T_662; 
  wire [63:0] _T_663; 
  wire  _T_665; 
  wire  _T_666; 
  wire  _T_667; 
  reg [4:0] _T_774; 
  reg [31:0] _RAND_13;
  wire  _T_775; 
  wire  _T_669; 
  wire [1:0] _T_777; 
  wire [2:0] _T_778; 
  wire [1:0] _T_779; 
  wire [1:0] _T_780; 
  wire [2:0] _T_782; 
  wire [1:0] _T_783; 
  wire [1:0] _T_784; 
  wire  _T_786; 
  reg  _T_818_1; 
  reg [31:0] _RAND_14;
  wire  _T_820_1; 
  wire  _T_822; 
  wire  _T_670; 
  wire [2:0] _GEN_0; 
  wire [2:0] _GEN_1; 
  wire [1:0] _T_703; 
  wire [3:0] _T_704; 
  wire [2:0] _T_705; 
  wire [2:0] _T_706; 
  wire  _T_707; 
  wire  _T_708; 
  wire  _T_709; 
  wire  _T_710; 
  wire  _T_712; 
  wire  _T_713; 
  wire  _T_715; 
  wire  _T_716; 
  wire  _T_717; 
  wire  _T_718; 
  wire  _T_719; 
  wire  _T_720; 
  wire  _T_721; 
  wire  _T_722; 
  wire  _T_723; 
  wire  _T_724; 
  wire  _T_725; 
  wire  _T_726; 
  wire  _T_727; 
  wire  _T_728; 
  wire  _T_729; 
  wire  _T_730; 
  wire  _T_731; 
  wire  _T_732; 
  wire  _T_733; 
  wire  _T_734; 
  wire  _T_735; 
  wire  _T_736; 
  wire  _T_737; 
  wire  _T_738; 
  wire  _T_739; 
  wire  _T_740; 
  wire  _T_741; 
  wire  _T_742; 
  wire  _T_743; 
  wire  _T_744; 
  wire  _T_745; 
  wire  _T_746; 
  wire  _T_747; 
  wire  _T_748; 
  wire  _T_749; 
  wire  _T_750; 
  wire  _T_751; 
  wire  _T_752; 
  wire  _T_753; 
  wire  _T_754; 
  wire  _T_755; 
  wire  _T_756; 
  wire  _T_757; 
  wire  _T_758; 
  wire [22:0] _T_767; 
  wire [7:0] _T_768; 
  wire [7:0] _T_769; 
  wire [4:0] _T_770; 
  wire  _T_771; 
  wire  _T_772; 
  wire  _T_776; 
  wire  _T_785; 
  wire  _T_788; 
  wire  _T_789; 
  wire  _T_792; 
  wire  _T_794; 
  wire  _T_797; 
  wire  _T_798; 
  wire  _T_801; 
  wire  _T_802; 
  wire  _T_803; 
  wire  _T_804; 
  wire  _T_806; 
  wire  _T_808; 
  wire  _T_809; 
  reg  _T_818_0; 
  reg [31:0] _RAND_15;
  wire  _T_824; 
  wire  _T_825; 
  wire  _T_826; 
  wire  _T_828; 
  wire  _T_813; 
  wire [4:0] _GEN_45; 
  wire [4:0] _T_815; 
  wire  _T_819_0; 
  wire  _T_819_1; 
  wire  _T_820_0; 
  wire  _T_821; 
  wire [64:0] _T_829; 
  wire [141:0] _T_832; 
  wire [190:0] _T_837; 
  wire [190:0] _T_838; 
  wire [190:0] _T_847; 
  wire [190:0] _T_848; 
  wire [190:0] _T_849; 
  wire  _T_862; 
  wire  _T_864; 
  wire [1:0] _T_865; 
  wire [2:0] _GEN_46; 
  wire  _T_866; 
  wire  _T_868; 
  wire  _T_870; 
  wire  _T_872; 
  wire  _T_874; 
  reg [4:0] _T_883; 
  reg [31:0] _RAND_16;
  wire  _T_886; 
  wire  _T_898; 
  wire  _T_904; 
  wire  _T_894; 
  wire  _T_895; 
  wire  _T_905; 
  wire  _T_910; 
  wire  _T_875; 
  wire [22:0] _T_877; 
  wire [7:0] _T_878; 
  wire [7:0] _T_879; 
  wire [4:0] _T_880; 
  wire  _T_881; 
  wire [4:0] _T_885; 
  wire  _T_899; 
  wire  _T_901; 
  wire  _T_902; 
  wire  _T_906; 
  wire  _T_907; 
  wire  _T_908; 
  wire  _T_911; 
  wire  _T_912; 
  dual_TLMonitor_14 dual_TLMonitor ( 
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_c_ready(TLMonitor_io_in_c_ready),
    .io_in_c_valid(TLMonitor_io_in_c_valid),
    .io_in_c_bits_opcode(TLMonitor_io_in_c_bits_opcode),
    .io_in_c_bits_param(TLMonitor_io_in_c_bits_param),
    .io_in_c_bits_size(TLMonitor_io_in_c_bits_size),
    .io_in_c_bits_source(TLMonitor_io_in_c_bits_source),
    .io_in_c_bits_address(TLMonitor_io_in_c_bits_address),
    .io_in_c_bits_corrupt(TLMonitor_io_in_c_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt),
    .io_in_e_ready(TLMonitor_io_in_e_ready),
    .io_in_e_valid(TLMonitor_io_in_e_valid),
    .io_in_e_bits_sink(TLMonitor_io_in_e_bits_sink)
  );
  assign _T_13 = _T_10_0_state == 2'h0; 
  assign _T_14 = _T_10_0_state == 2'h2; 
  assign _T_15 = _T_10_0_state == 2'h3; 
  assign _T_17 = _T_15 | _T_14; 
  assign _T_18 = _T_10_0_state != 2'h0; 
  assign _T_25 = auto_in_a_bits_address ^ 32'h40000000; 
  assign _T_26 = {1'b0,$signed(_T_25)}; 
  assign _T_27 = $signed(_T_26) & $signed(33'shc0000000); 
  assign _T_28 = $signed(_T_27); 
  assign _T_29 = $signed(_T_28) == $signed(33'sh0); 
  assign _T_37 = {1'b0,$signed(auto_in_a_bits_address)}; 
  assign _T_38 = $signed(_T_37) & $signed(33'shc0000000); 
  assign _T_39 = $signed(_T_38); 
  assign _T_40 = $signed(_T_39) == $signed(33'sh0); 
  assign _T_71 = auto_in_a_bits_opcode == 3'h3; 
  assign _T_72 = auto_in_a_bits_opcode == 3'h2; 
  assign _T_73 = _T_72 ? 1'h0 : 1'h1; 
  assign _T_74 = _T_71 ? 1'h0 : _T_73; 
  assign _T_95 = _T_40 ? 2'h2 : 2'h0; 
  assign _GEN_43 = {{1'd0}, _T_29}; 
  assign _T_97 = _GEN_43 | _T_95; 
  assign _T_99 = _T_11_0_fifoId == _T_97; 
  assign _T_100 = _T_17 & _T_99; 
  assign _T_104 = _T_11_0_bits_data[0]; 
  assign _T_105 = _T_12_0_data[0]; 
  assign _T_106 = {_T_104,_T_105}; 
  assign _T_107 = _T_11_0_bits_data[1]; 
  assign _T_108 = _T_12_0_data[1]; 
  assign _T_109 = {_T_107,_T_108}; 
  assign _T_110 = _T_11_0_bits_data[2]; 
  assign _T_111 = _T_12_0_data[2]; 
  assign _T_112 = {_T_110,_T_111}; 
  assign _T_113 = _T_11_0_bits_data[3]; 
  assign _T_114 = _T_12_0_data[3]; 
  assign _T_115 = {_T_113,_T_114}; 
  assign _T_116 = _T_11_0_bits_data[4]; 
  assign _T_117 = _T_12_0_data[4]; 
  assign _T_118 = {_T_116,_T_117}; 
  assign _T_119 = _T_11_0_bits_data[5]; 
  assign _T_120 = _T_12_0_data[5]; 
  assign _T_121 = {_T_119,_T_120}; 
  assign _T_122 = _T_11_0_bits_data[6]; 
  assign _T_123 = _T_12_0_data[6]; 
  assign _T_124 = {_T_122,_T_123}; 
  assign _T_125 = _T_11_0_bits_data[7]; 
  assign _T_126 = _T_12_0_data[7]; 
  assign _T_127 = {_T_125,_T_126}; 
  assign _T_128 = _T_11_0_bits_data[8]; 
  assign _T_129 = _T_12_0_data[8]; 
  assign _T_130 = {_T_128,_T_129}; 
  assign _T_131 = _T_11_0_bits_data[9]; 
  assign _T_132 = _T_12_0_data[9]; 
  assign _T_133 = {_T_131,_T_132}; 
  assign _T_134 = _T_11_0_bits_data[10]; 
  assign _T_135 = _T_12_0_data[10]; 
  assign _T_136 = {_T_134,_T_135}; 
  assign _T_137 = _T_11_0_bits_data[11]; 
  assign _T_138 = _T_12_0_data[11]; 
  assign _T_139 = {_T_137,_T_138}; 
  assign _T_140 = _T_11_0_bits_data[12]; 
  assign _T_141 = _T_12_0_data[12]; 
  assign _T_142 = {_T_140,_T_141}; 
  assign _T_143 = _T_11_0_bits_data[13]; 
  assign _T_144 = _T_12_0_data[13]; 
  assign _T_145 = {_T_143,_T_144}; 
  assign _T_146 = _T_11_0_bits_data[14]; 
  assign _T_147 = _T_12_0_data[14]; 
  assign _T_148 = {_T_146,_T_147}; 
  assign _T_149 = _T_11_0_bits_data[15]; 
  assign _T_150 = _T_12_0_data[15]; 
  assign _T_151 = {_T_149,_T_150}; 
  assign _T_152 = _T_11_0_bits_data[16]; 
  assign _T_153 = _T_12_0_data[16]; 
  assign _T_154 = {_T_152,_T_153}; 
  assign _T_155 = _T_11_0_bits_data[17]; 
  assign _T_156 = _T_12_0_data[17]; 
  assign _T_157 = {_T_155,_T_156}; 
  assign _T_158 = _T_11_0_bits_data[18]; 
  assign _T_159 = _T_12_0_data[18]; 
  assign _T_160 = {_T_158,_T_159}; 
  assign _T_161 = _T_11_0_bits_data[19]; 
  assign _T_162 = _T_12_0_data[19]; 
  assign _T_163 = {_T_161,_T_162}; 
  assign _T_164 = _T_11_0_bits_data[20]; 
  assign _T_165 = _T_12_0_data[20]; 
  assign _T_166 = {_T_164,_T_165}; 
  assign _T_167 = _T_11_0_bits_data[21]; 
  assign _T_168 = _T_12_0_data[21]; 
  assign _T_169 = {_T_167,_T_168}; 
  assign _T_170 = _T_11_0_bits_data[22]; 
  assign _T_171 = _T_12_0_data[22]; 
  assign _T_172 = {_T_170,_T_171}; 
  assign _T_173 = _T_11_0_bits_data[23]; 
  assign _T_174 = _T_12_0_data[23]; 
  assign _T_175 = {_T_173,_T_174}; 
  assign _T_176 = _T_11_0_bits_data[24]; 
  assign _T_177 = _T_12_0_data[24]; 
  assign _T_178 = {_T_176,_T_177}; 
  assign _T_179 = _T_11_0_bits_data[25]; 
  assign _T_180 = _T_12_0_data[25]; 
  assign _T_181 = {_T_179,_T_180}; 
  assign _T_182 = _T_11_0_bits_data[26]; 
  assign _T_183 = _T_12_0_data[26]; 
  assign _T_184 = {_T_182,_T_183}; 
  assign _T_185 = _T_11_0_bits_data[27]; 
  assign _T_186 = _T_12_0_data[27]; 
  assign _T_187 = {_T_185,_T_186}; 
  assign _T_188 = _T_11_0_bits_data[28]; 
  assign _T_189 = _T_12_0_data[28]; 
  assign _T_190 = {_T_188,_T_189}; 
  assign _T_191 = _T_11_0_bits_data[29]; 
  assign _T_192 = _T_12_0_data[29]; 
  assign _T_193 = {_T_191,_T_192}; 
  assign _T_194 = _T_11_0_bits_data[30]; 
  assign _T_195 = _T_12_0_data[30]; 
  assign _T_196 = {_T_194,_T_195}; 
  assign _T_197 = _T_11_0_bits_data[31]; 
  assign _T_198 = _T_12_0_data[31]; 
  assign _T_199 = {_T_197,_T_198}; 
  assign _T_200 = _T_11_0_bits_data[32]; 
  assign _T_201 = _T_12_0_data[32]; 
  assign _T_202 = {_T_200,_T_201}; 
  assign _T_203 = _T_11_0_bits_data[33]; 
  assign _T_204 = _T_12_0_data[33]; 
  assign _T_205 = {_T_203,_T_204}; 
  assign _T_206 = _T_11_0_bits_data[34]; 
  assign _T_207 = _T_12_0_data[34]; 
  assign _T_208 = {_T_206,_T_207}; 
  assign _T_209 = _T_11_0_bits_data[35]; 
  assign _T_210 = _T_12_0_data[35]; 
  assign _T_211 = {_T_209,_T_210}; 
  assign _T_212 = _T_11_0_bits_data[36]; 
  assign _T_213 = _T_12_0_data[36]; 
  assign _T_214 = {_T_212,_T_213}; 
  assign _T_215 = _T_11_0_bits_data[37]; 
  assign _T_216 = _T_12_0_data[37]; 
  assign _T_217 = {_T_215,_T_216}; 
  assign _T_218 = _T_11_0_bits_data[38]; 
  assign _T_219 = _T_12_0_data[38]; 
  assign _T_220 = {_T_218,_T_219}; 
  assign _T_221 = _T_11_0_bits_data[39]; 
  assign _T_222 = _T_12_0_data[39]; 
  assign _T_223 = {_T_221,_T_222}; 
  assign _T_224 = _T_11_0_bits_data[40]; 
  assign _T_225 = _T_12_0_data[40]; 
  assign _T_226 = {_T_224,_T_225}; 
  assign _T_227 = _T_11_0_bits_data[41]; 
  assign _T_228 = _T_12_0_data[41]; 
  assign _T_229 = {_T_227,_T_228}; 
  assign _T_230 = _T_11_0_bits_data[42]; 
  assign _T_231 = _T_12_0_data[42]; 
  assign _T_232 = {_T_230,_T_231}; 
  assign _T_233 = _T_11_0_bits_data[43]; 
  assign _T_234 = _T_12_0_data[43]; 
  assign _T_235 = {_T_233,_T_234}; 
  assign _T_236 = _T_11_0_bits_data[44]; 
  assign _T_237 = _T_12_0_data[44]; 
  assign _T_238 = {_T_236,_T_237}; 
  assign _T_239 = _T_11_0_bits_data[45]; 
  assign _T_240 = _T_12_0_data[45]; 
  assign _T_241 = {_T_239,_T_240}; 
  assign _T_242 = _T_11_0_bits_data[46]; 
  assign _T_243 = _T_12_0_data[46]; 
  assign _T_244 = {_T_242,_T_243}; 
  assign _T_245 = _T_11_0_bits_data[47]; 
  assign _T_246 = _T_12_0_data[47]; 
  assign _T_247 = {_T_245,_T_246}; 
  assign _T_248 = _T_11_0_bits_data[48]; 
  assign _T_249 = _T_12_0_data[48]; 
  assign _T_250 = {_T_248,_T_249}; 
  assign _T_251 = _T_11_0_bits_data[49]; 
  assign _T_252 = _T_12_0_data[49]; 
  assign _T_253 = {_T_251,_T_252}; 
  assign _T_254 = _T_11_0_bits_data[50]; 
  assign _T_255 = _T_12_0_data[50]; 
  assign _T_256 = {_T_254,_T_255}; 
  assign _T_257 = _T_11_0_bits_data[51]; 
  assign _T_258 = _T_12_0_data[51]; 
  assign _T_259 = {_T_257,_T_258}; 
  assign _T_260 = _T_11_0_bits_data[52]; 
  assign _T_261 = _T_12_0_data[52]; 
  assign _T_262 = {_T_260,_T_261}; 
  assign _T_263 = _T_11_0_bits_data[53]; 
  assign _T_264 = _T_12_0_data[53]; 
  assign _T_265 = {_T_263,_T_264}; 
  assign _T_266 = _T_11_0_bits_data[54]; 
  assign _T_267 = _T_12_0_data[54]; 
  assign _T_268 = {_T_266,_T_267}; 
  assign _T_269 = _T_11_0_bits_data[55]; 
  assign _T_270 = _T_12_0_data[55]; 
  assign _T_271 = {_T_269,_T_270}; 
  assign _T_272 = _T_11_0_bits_data[56]; 
  assign _T_273 = _T_12_0_data[56]; 
  assign _T_274 = {_T_272,_T_273}; 
  assign _T_275 = _T_11_0_bits_data[57]; 
  assign _T_276 = _T_12_0_data[57]; 
  assign _T_277 = {_T_275,_T_276}; 
  assign _T_278 = _T_11_0_bits_data[58]; 
  assign _T_279 = _T_12_0_data[58]; 
  assign _T_280 = {_T_278,_T_279}; 
  assign _T_281 = _T_11_0_bits_data[59]; 
  assign _T_282 = _T_12_0_data[59]; 
  assign _T_283 = {_T_281,_T_282}; 
  assign _T_284 = _T_11_0_bits_data[60]; 
  assign _T_285 = _T_12_0_data[60]; 
  assign _T_286 = {_T_284,_T_285}; 
  assign _T_287 = _T_11_0_bits_data[61]; 
  assign _T_288 = _T_12_0_data[61]; 
  assign _T_289 = {_T_287,_T_288}; 
  assign _T_290 = _T_11_0_bits_data[62]; 
  assign _T_291 = _T_12_0_data[62]; 
  assign _T_292 = {_T_290,_T_291}; 
  assign _T_293 = _T_11_0_bits_data[63]; 
  assign _T_294 = _T_12_0_data[63]; 
  assign _T_295 = {_T_293,_T_294}; 
  assign _T_296 = _T_11_0_lut >> _T_106; 
  assign _T_297 = _T_296[0]; 
  assign _T_298 = _T_11_0_lut >> _T_109; 
  assign _T_299 = _T_298[0]; 
  assign _T_300 = _T_11_0_lut >> _T_112; 
  assign _T_301 = _T_300[0]; 
  assign _T_302 = _T_11_0_lut >> _T_115; 
  assign _T_303 = _T_302[0]; 
  assign _T_304 = _T_11_0_lut >> _T_118; 
  assign _T_305 = _T_304[0]; 
  assign _T_306 = _T_11_0_lut >> _T_121; 
  assign _T_307 = _T_306[0]; 
  assign _T_308 = _T_11_0_lut >> _T_124; 
  assign _T_309 = _T_308[0]; 
  assign _T_310 = _T_11_0_lut >> _T_127; 
  assign _T_311 = _T_310[0]; 
  assign _T_312 = _T_11_0_lut >> _T_130; 
  assign _T_313 = _T_312[0]; 
  assign _T_314 = _T_11_0_lut >> _T_133; 
  assign _T_315 = _T_314[0]; 
  assign _T_316 = _T_11_0_lut >> _T_136; 
  assign _T_317 = _T_316[0]; 
  assign _T_318 = _T_11_0_lut >> _T_139; 
  assign _T_319 = _T_318[0]; 
  assign _T_320 = _T_11_0_lut >> _T_142; 
  assign _T_321 = _T_320[0]; 
  assign _T_322 = _T_11_0_lut >> _T_145; 
  assign _T_323 = _T_322[0]; 
  assign _T_324 = _T_11_0_lut >> _T_148; 
  assign _T_325 = _T_324[0]; 
  assign _T_326 = _T_11_0_lut >> _T_151; 
  assign _T_327 = _T_326[0]; 
  assign _T_328 = _T_11_0_lut >> _T_154; 
  assign _T_329 = _T_328[0]; 
  assign _T_330 = _T_11_0_lut >> _T_157; 
  assign _T_331 = _T_330[0]; 
  assign _T_332 = _T_11_0_lut >> _T_160; 
  assign _T_333 = _T_332[0]; 
  assign _T_334 = _T_11_0_lut >> _T_163; 
  assign _T_335 = _T_334[0]; 
  assign _T_336 = _T_11_0_lut >> _T_166; 
  assign _T_337 = _T_336[0]; 
  assign _T_338 = _T_11_0_lut >> _T_169; 
  assign _T_339 = _T_338[0]; 
  assign _T_340 = _T_11_0_lut >> _T_172; 
  assign _T_341 = _T_340[0]; 
  assign _T_342 = _T_11_0_lut >> _T_175; 
  assign _T_343 = _T_342[0]; 
  assign _T_344 = _T_11_0_lut >> _T_178; 
  assign _T_345 = _T_344[0]; 
  assign _T_346 = _T_11_0_lut >> _T_181; 
  assign _T_347 = _T_346[0]; 
  assign _T_348 = _T_11_0_lut >> _T_184; 
  assign _T_349 = _T_348[0]; 
  assign _T_350 = _T_11_0_lut >> _T_187; 
  assign _T_351 = _T_350[0]; 
  assign _T_352 = _T_11_0_lut >> _T_190; 
  assign _T_353 = _T_352[0]; 
  assign _T_354 = _T_11_0_lut >> _T_193; 
  assign _T_355 = _T_354[0]; 
  assign _T_356 = _T_11_0_lut >> _T_196; 
  assign _T_357 = _T_356[0]; 
  assign _T_358 = _T_11_0_lut >> _T_199; 
  assign _T_359 = _T_358[0]; 
  assign _T_360 = _T_11_0_lut >> _T_202; 
  assign _T_361 = _T_360[0]; 
  assign _T_362 = _T_11_0_lut >> _T_205; 
  assign _T_363 = _T_362[0]; 
  assign _T_364 = _T_11_0_lut >> _T_208; 
  assign _T_365 = _T_364[0]; 
  assign _T_366 = _T_11_0_lut >> _T_211; 
  assign _T_367 = _T_366[0]; 
  assign _T_368 = _T_11_0_lut >> _T_214; 
  assign _T_369 = _T_368[0]; 
  assign _T_370 = _T_11_0_lut >> _T_217; 
  assign _T_371 = _T_370[0]; 
  assign _T_372 = _T_11_0_lut >> _T_220; 
  assign _T_373 = _T_372[0]; 
  assign _T_374 = _T_11_0_lut >> _T_223; 
  assign _T_375 = _T_374[0]; 
  assign _T_376 = _T_11_0_lut >> _T_226; 
  assign _T_377 = _T_376[0]; 
  assign _T_378 = _T_11_0_lut >> _T_229; 
  assign _T_379 = _T_378[0]; 
  assign _T_380 = _T_11_0_lut >> _T_232; 
  assign _T_381 = _T_380[0]; 
  assign _T_382 = _T_11_0_lut >> _T_235; 
  assign _T_383 = _T_382[0]; 
  assign _T_384 = _T_11_0_lut >> _T_238; 
  assign _T_385 = _T_384[0]; 
  assign _T_386 = _T_11_0_lut >> _T_241; 
  assign _T_387 = _T_386[0]; 
  assign _T_388 = _T_11_0_lut >> _T_244; 
  assign _T_389 = _T_388[0]; 
  assign _T_390 = _T_11_0_lut >> _T_247; 
  assign _T_391 = _T_390[0]; 
  assign _T_392 = _T_11_0_lut >> _T_250; 
  assign _T_393 = _T_392[0]; 
  assign _T_394 = _T_11_0_lut >> _T_253; 
  assign _T_395 = _T_394[0]; 
  assign _T_396 = _T_11_0_lut >> _T_256; 
  assign _T_397 = _T_396[0]; 
  assign _T_398 = _T_11_0_lut >> _T_259; 
  assign _T_399 = _T_398[0]; 
  assign _T_400 = _T_11_0_lut >> _T_262; 
  assign _T_401 = _T_400[0]; 
  assign _T_402 = _T_11_0_lut >> _T_265; 
  assign _T_403 = _T_402[0]; 
  assign _T_404 = _T_11_0_lut >> _T_268; 
  assign _T_405 = _T_404[0]; 
  assign _T_406 = _T_11_0_lut >> _T_271; 
  assign _T_407 = _T_406[0]; 
  assign _T_408 = _T_11_0_lut >> _T_274; 
  assign _T_409 = _T_408[0]; 
  assign _T_410 = _T_11_0_lut >> _T_277; 
  assign _T_411 = _T_410[0]; 
  assign _T_412 = _T_11_0_lut >> _T_280; 
  assign _T_413 = _T_412[0]; 
  assign _T_414 = _T_11_0_lut >> _T_283; 
  assign _T_415 = _T_414[0]; 
  assign _T_416 = _T_11_0_lut >> _T_286; 
  assign _T_417 = _T_416[0]; 
  assign _T_418 = _T_11_0_lut >> _T_289; 
  assign _T_419 = _T_418[0]; 
  assign _T_420 = _T_11_0_lut >> _T_292; 
  assign _T_421 = _T_420[0]; 
  assign _T_422 = _T_11_0_lut >> _T_295; 
  assign _T_423 = _T_422[0]; 
  assign _T_430 = {_T_311,_T_309,_T_307,_T_305,_T_303,_T_301,_T_299,_T_297}; 
  assign _T_438 = {_T_327,_T_325,_T_323,_T_321,_T_319,_T_317,_T_315,_T_313,_T_430}; 
  assign _T_445 = {_T_343,_T_341,_T_339,_T_337,_T_335,_T_333,_T_331,_T_329}; 
  assign _T_454 = {_T_359,_T_357,_T_355,_T_353,_T_351,_T_349,_T_347,_T_345,_T_445,_T_438}; 
  assign _T_461 = {_T_375,_T_373,_T_371,_T_369,_T_367,_T_365,_T_363,_T_361}; 
  assign _T_469 = {_T_391,_T_389,_T_387,_T_385,_T_383,_T_381,_T_379,_T_377,_T_461}; 
  assign _T_476 = {_T_407,_T_405,_T_403,_T_401,_T_399,_T_397,_T_395,_T_393}; 
  assign _T_485 = {_T_423,_T_421,_T_419,_T_417,_T_415,_T_413,_T_411,_T_409,_T_476,_T_469}; 
  assign _T_486 = {_T_485,_T_454}; 
  assign _T_487 = _T_11_0_bits_param[1]; 
  assign _T_488 = _T_11_0_bits_param[0]; 
  assign _T_489 = _T_11_0_bits_param[2]; 
  assign _T_490 = ~ _T_11_0_bits_mask; 
  assign _T_491 = _T_11_0_bits_mask[7:1]; 
  assign _GEN_44 = {{1'd0}, _T_491}; 
  assign _T_492 = _T_490 | _GEN_44; 
  assign _T_493 = ~ _T_492; 
  assign _T_508 = {_T_293,_T_269,_T_245,_T_221,_T_197,_T_173,_T_149,_T_125}; 
  assign _T_523 = {_T_294,_T_270,_T_246,_T_222,_T_198,_T_174,_T_150,_T_126}; 
  assign _T_524 = _T_508 & _T_493; 
  assign _T_525 = {_T_524, 1'h0}; 
  assign _T_526 = _T_525[7:0]; 
  assign _T_527 = _T_523 & _T_493; 
  assign _T_528 = {_T_527, 1'h0}; 
  assign _T_529 = _T_528[7:0]; 
  assign _T_530 = {_T_526, 1'h0}; 
  assign _T_531 = _T_530[7:0]; 
  assign _T_532 = _T_526 | _T_531; 
  assign _T_533 = {_T_532, 2'h0}; 
  assign _T_534 = _T_533[7:0]; 
  assign _T_535 = _T_532 | _T_534; 
  assign _T_536 = {_T_535, 4'h0}; 
  assign _T_537 = _T_536[7:0]; 
  assign _T_538 = _T_535 | _T_537; 
  assign _T_540 = _T_538[0]; 
  assign _T_541 = _T_538[1]; 
  assign _T_542 = _T_538[2]; 
  assign _T_543 = _T_538[3]; 
  assign _T_544 = _T_538[4]; 
  assign _T_545 = _T_538[5]; 
  assign _T_546 = _T_538[6]; 
  assign _T_547 = _T_538[7]; 
  assign _T_549 = _T_540 ? 8'hff : 8'h0; 
  assign _T_551 = _T_541 ? 8'hff : 8'h0; 
  assign _T_553 = _T_542 ? 8'hff : 8'h0; 
  assign _T_555 = _T_543 ? 8'hff : 8'h0; 
  assign _T_557 = _T_544 ? 8'hff : 8'h0; 
  assign _T_559 = _T_545 ? 8'hff : 8'h0; 
  assign _T_561 = _T_546 ? 8'hff : 8'h0; 
  assign _T_563 = _T_547 ? 8'hff : 8'h0; 
  assign _T_570 = {_T_563,_T_561,_T_559,_T_557,_T_555,_T_553,_T_551,_T_549}; 
  assign _T_571 = {_T_529, 1'h0}; 
  assign _T_572 = _T_571[7:0]; 
  assign _T_573 = _T_529 | _T_572; 
  assign _T_574 = {_T_573, 2'h0}; 
  assign _T_575 = _T_574[7:0]; 
  assign _T_576 = _T_573 | _T_575; 
  assign _T_577 = {_T_576, 4'h0}; 
  assign _T_578 = _T_577[7:0]; 
  assign _T_579 = _T_576 | _T_578; 
  assign _T_581 = _T_579[0]; 
  assign _T_582 = _T_579[1]; 
  assign _T_583 = _T_579[2]; 
  assign _T_584 = _T_579[3]; 
  assign _T_585 = _T_579[4]; 
  assign _T_586 = _T_579[5]; 
  assign _T_587 = _T_579[6]; 
  assign _T_588 = _T_579[7]; 
  assign _T_590 = _T_581 ? 8'hff : 8'h0; 
  assign _T_592 = _T_582 ? 8'hff : 8'h0; 
  assign _T_594 = _T_583 ? 8'hff : 8'h0; 
  assign _T_596 = _T_584 ? 8'hff : 8'h0; 
  assign _T_598 = _T_585 ? 8'hff : 8'h0; 
  assign _T_600 = _T_586 ? 8'hff : 8'h0; 
  assign _T_602 = _T_587 ? 8'hff : 8'h0; 
  assign _T_604 = _T_588 ? 8'hff : 8'h0; 
  assign _T_611 = {_T_604,_T_602,_T_600,_T_598,_T_596,_T_594,_T_592,_T_590}; 
  assign _T_612 = _T_11_0_bits_mask[0]; 
  assign _T_613 = _T_11_0_bits_mask[1]; 
  assign _T_614 = _T_11_0_bits_mask[2]; 
  assign _T_615 = _T_11_0_bits_mask[3]; 
  assign _T_616 = _T_11_0_bits_mask[4]; 
  assign _T_617 = _T_11_0_bits_mask[5]; 
  assign _T_618 = _T_11_0_bits_mask[6]; 
  assign _T_619 = _T_11_0_bits_mask[7]; 
  assign _T_621 = _T_612 ? 8'hff : 8'h0; 
  assign _T_623 = _T_613 ? 8'hff : 8'h0; 
  assign _T_625 = _T_614 ? 8'hff : 8'h0; 
  assign _T_627 = _T_615 ? 8'hff : 8'h0; 
  assign _T_629 = _T_616 ? 8'hff : 8'h0; 
  assign _T_631 = _T_617 ? 8'hff : 8'h0; 
  assign _T_633 = _T_618 ? 8'hff : 8'h0; 
  assign _T_635 = _T_619 ? 8'hff : 8'h0; 
  assign _T_642 = {_T_635,_T_633,_T_631,_T_629,_T_627,_T_625,_T_623,_T_621}; 
  assign _T_643 = _T_11_0_bits_data & _T_642; 
  assign _T_644 = _T_643 | _T_570; 
  assign _T_645 = _T_12_0_data & _T_642; 
  assign _T_646 = _T_645 | _T_611; 
  assign _T_647 = ~ _T_646; 
  assign _T_648 = _T_489 ? _T_646 : _T_647; 
  assign _T_650 = _T_644 + _T_648; 
  assign _T_651 = _T_644[63]; 
  assign _T_652 = _T_487 == _T_651; 
  assign _T_654 = _T_646[63]; 
  assign _T_655 = _T_651 == _T_654; 
  assign _T_656 = _T_650[63]; 
  assign _T_657 = _T_656 == 1'h0; 
  assign _T_658 = _T_655 ? _T_657 : _T_652; 
  assign _T_659 = _T_488 == _T_658; 
  assign _T_660 = _T_659 ? _T_11_0_bits_data : _T_12_0_data; 
  assign _T_661 = _T_489 ? _T_650 : _T_660; 
  assign _T_662 = _T_11_0_bits_opcode[0]; 
  assign _T_663 = _T_662 ? _T_486 : _T_661; 
  assign _T_665 = _T_100 == 1'h0; 
  assign _T_666 = _T_74 | _T_13; 
  assign _T_667 = _T_665 & _T_666; 
  assign _T_775 = _T_774 == 5'h0; 
  assign _T_669 = auto_in_a_valid & _T_667; 
  assign _T_777 = {_T_669,_T_14}; 
  assign _T_778 = {_T_777, 1'h0}; 
  assign _T_779 = _T_778[1:0]; 
  assign _T_780 = _T_777 | _T_779; 
  assign _T_782 = {_T_780, 1'h0}; 
  assign _T_783 = _T_782[1:0]; 
  assign _T_784 = ~ _T_783; 
  assign _T_786 = _T_784[1]; 
  assign _T_820_1 = _T_775 ? _T_786 : _T_818_1; 
  assign _T_822 = auto_out_a_ready & _T_820_1; 
  assign _T_670 = _T_74 == 1'h0; 
  assign _GEN_0 = _T_670 ? 3'h4 : auto_in_a_bits_opcode; 
  assign _GEN_1 = _T_670 ? 3'h0 : auto_in_a_bits_param; 
  assign _T_703 = _T_11_0_bits_size[1:0]; 
  assign _T_704 = 4'h1 << _T_703; 
  assign _T_705 = _T_704[2:0]; 
  assign _T_706 = _T_705 | 3'h1; 
  assign _T_707 = _T_11_0_bits_size >= 4'h3; 
  assign _T_708 = _T_706[2]; 
  assign _T_709 = _T_11_0_bits_address[2]; 
  assign _T_710 = _T_709 == 1'h0; 
  assign _T_712 = _T_708 & _T_710; 
  assign _T_713 = _T_707 | _T_712; 
  assign _T_715 = _T_708 & _T_709; 
  assign _T_716 = _T_707 | _T_715; 
  assign _T_717 = _T_706[1]; 
  assign _T_718 = _T_11_0_bits_address[1]; 
  assign _T_719 = _T_718 == 1'h0; 
  assign _T_720 = _T_710 & _T_719; 
  assign _T_721 = _T_717 & _T_720; 
  assign _T_722 = _T_713 | _T_721; 
  assign _T_723 = _T_710 & _T_718; 
  assign _T_724 = _T_717 & _T_723; 
  assign _T_725 = _T_713 | _T_724; 
  assign _T_726 = _T_709 & _T_719; 
  assign _T_727 = _T_717 & _T_726; 
  assign _T_728 = _T_716 | _T_727; 
  assign _T_729 = _T_709 & _T_718; 
  assign _T_730 = _T_717 & _T_729; 
  assign _T_731 = _T_716 | _T_730; 
  assign _T_732 = _T_706[0]; 
  assign _T_733 = _T_11_0_bits_address[0]; 
  assign _T_734 = _T_733 == 1'h0; 
  assign _T_735 = _T_720 & _T_734; 
  assign _T_736 = _T_732 & _T_735; 
  assign _T_737 = _T_722 | _T_736; 
  assign _T_738 = _T_720 & _T_733; 
  assign _T_739 = _T_732 & _T_738; 
  assign _T_740 = _T_722 | _T_739; 
  assign _T_741 = _T_723 & _T_734; 
  assign _T_742 = _T_732 & _T_741; 
  assign _T_743 = _T_725 | _T_742; 
  assign _T_744 = _T_723 & _T_733; 
  assign _T_745 = _T_732 & _T_744; 
  assign _T_746 = _T_725 | _T_745; 
  assign _T_747 = _T_726 & _T_734; 
  assign _T_748 = _T_732 & _T_747; 
  assign _T_749 = _T_728 | _T_748; 
  assign _T_750 = _T_726 & _T_733; 
  assign _T_751 = _T_732 & _T_750; 
  assign _T_752 = _T_728 | _T_751; 
  assign _T_753 = _T_729 & _T_734; 
  assign _T_754 = _T_732 & _T_753; 
  assign _T_755 = _T_731 | _T_754; 
  assign _T_756 = _T_729 & _T_733; 
  assign _T_757 = _T_732 & _T_756; 
  assign _T_758 = _T_731 | _T_757; 
  assign _T_767 = 23'hff << auto_in_a_bits_size; 
  assign _T_768 = _T_767[7:0]; 
  assign _T_769 = ~ _T_768; 
  assign _T_770 = _T_769[7:3]; 
  assign _T_771 = auto_in_a_bits_opcode[2]; 
  assign _T_772 = _T_771 == 1'h0; 
  assign _T_776 = _T_775 & auto_out_a_ready; 
  assign _T_785 = _T_784[0]; 
  assign _T_788 = _T_785 & _T_14; 
  assign _T_789 = _T_786 & _T_669; 
  assign _T_792 = _T_788 | _T_789; 
  assign _T_794 = _T_788 == 1'h0; 
  assign _T_797 = _T_789 == 1'h0; 
  assign _T_798 = _T_794 | _T_797; 
  assign _T_801 = _T_798 | reset; 
  assign _T_802 = _T_801 == 1'h0; 
  assign _T_803 = _T_14 | _T_669; 
  assign _T_804 = _T_803 == 1'h0; 
  assign _T_806 = _T_804 | _T_792; 
  assign _T_808 = _T_806 | reset; 
  assign _T_809 = _T_808 == 1'h0; 
  assign _T_824 = _T_818_0 ? _T_14 : 1'h0; 
  assign _T_825 = _T_818_1 ? _T_669 : 1'h0; 
  assign _T_826 = _T_824 | _T_825; 
  assign _T_828 = _T_775 ? _T_803 : _T_826; 
  assign _T_813 = auto_out_a_ready & _T_828; 
  assign _GEN_45 = {{4'd0}, _T_813}; 
  assign _T_815 = _T_774 - _GEN_45; 
  assign _T_819_0 = _T_775 ? _T_788 : _T_818_0; 
  assign _T_819_1 = _T_775 ? _T_789 : _T_818_1; 
  assign _T_820_0 = _T_775 ? _T_785 : _T_818_0; 
  assign _T_821 = auto_out_a_ready & _T_820_0; 
  assign _T_829 = {_T_663,_T_12_0_corrupt}; 
  assign _T_832 = {69'h0,_T_758,_T_755,_T_752,_T_749,_T_746,_T_743,_T_740,_T_737,_T_829}; 
  assign _T_837 = {6'h0,_T_11_0_bits_size,_T_11_0_bits_source,_T_11_0_bits_address,_T_832}; 
  assign _T_838 = _T_819_0 ? _T_837 : 191'h0; 
  assign _T_847 = {_GEN_0,_GEN_1,auto_in_a_bits_size,auto_in_a_bits_source,auto_in_a_bits_address,69'h0,auto_in_a_bits_mask,auto_in_a_bits_data,1'h0}; 
  assign _T_848 = _T_819_1 ? _T_847 : 191'h0; 
  assign _T_849 = _T_838 | _T_848; 
  assign _T_862 = _T_822 & _T_669; 
  assign _T_864 = _T_862 & _T_670; 
  assign _T_865 = auto_in_a_bits_param[1:0]; 
  assign _GEN_46 = {{1'd0}, _T_865}; 
  assign _T_866 = 3'h3 == _GEN_46; 
  assign _T_868 = 3'h0 == _GEN_46; 
  assign _T_870 = 3'h1 == _GEN_46; 
  assign _T_872 = 3'h2 == _GEN_46; 
  assign _T_874 = _T_821 & _T_14; 
  assign _T_886 = _T_883 == 5'h0; 
  assign _T_898 = auto_out_d_bits_opcode == 3'h1; 
  assign _T_904 = _T_886 & _T_898; 
  assign _T_894 = _T_11_0_bits_source == auto_out_d_bits_source; 
  assign _T_895 = _T_894 & _T_18; 
  assign _T_905 = _T_904 & _T_895; 
  assign _T_910 = auto_in_d_ready | _T_905; 
  assign _T_875 = _T_910 & auto_out_d_valid; 
  assign _T_877 = 23'hff << auto_out_d_bits_size; 
  assign _T_878 = _T_877[7:0]; 
  assign _T_879 = ~ _T_878; 
  assign _T_880 = _T_879[7:3]; 
  assign _T_881 = auto_out_d_bits_opcode[0]; 
  assign _T_885 = _T_883 - 5'h1; 
  assign _T_899 = auto_out_d_bits_opcode == 3'h0; 
  assign _T_901 = _T_875 & _T_886; 
  assign _T_902 = _T_895 & _T_898; 
  assign _T_906 = _T_886 & _T_899; 
  assign _T_907 = _T_906 & _T_895; 
  assign _T_908 = _T_905 == 1'h0; 
  assign _T_911 = _T_12_0_corrupt | auto_out_d_bits_denied; 
  assign _T_912 = _T_12_0_denied | auto_out_d_bits_denied; 
  assign auto_in_a_ready = _T_822 & _T_667; 
  assign auto_in_c_ready = auto_out_c_ready; 
  assign auto_in_d_valid = auto_out_d_valid & _T_908; 
  assign auto_in_d_bits_opcode = _T_907 ? 3'h1 : auto_out_d_bits_opcode; 
  assign auto_in_d_bits_param = auto_out_d_bits_param; 
  assign auto_in_d_bits_size = auto_out_d_bits_size; 
  assign auto_in_d_bits_source = auto_out_d_bits_source; 
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; 
  assign auto_in_d_bits_denied = _T_907 ? _T_912 : auto_out_d_bits_denied; 
  assign auto_in_d_bits_data = _T_907 ? _T_12_0_data : auto_out_d_bits_data; 
  assign auto_in_d_bits_corrupt = _T_907 ? _T_911 : auto_out_d_bits_corrupt; 
  assign auto_in_e_ready = auto_out_e_ready; 
  assign auto_out_a_valid = _T_775 ? _T_803 : _T_826; 
  assign auto_out_a_bits_opcode = _T_849[190:188]; 
  assign auto_out_a_bits_param = _T_849[187:185]; 
  assign auto_out_a_bits_size = _T_849[184:181]; 
  assign auto_out_a_bits_source = _T_849[180:174]; 
  assign auto_out_a_bits_address = _T_849[173:142]; 
  assign auto_out_a_bits_mask = _T_849[72:65]; 
  assign auto_out_a_bits_data = _T_849[64:1]; 
  assign auto_out_a_bits_corrupt = _T_849[0]; 
  assign auto_out_c_valid = auto_in_c_valid; 
  assign auto_out_c_bits_opcode = auto_in_c_bits_opcode; 
  assign auto_out_c_bits_param = auto_in_c_bits_param; 
  assign auto_out_c_bits_size = auto_in_c_bits_size; 
  assign auto_out_c_bits_source = auto_in_c_bits_source; 
  assign auto_out_c_bits_address = auto_in_c_bits_address; 
  assign auto_out_c_bits_corrupt = auto_in_c_bits_corrupt; 
  assign auto_out_d_ready = auto_in_d_ready | _T_905; 
  assign auto_out_e_valid = auto_in_e_valid; 
  assign auto_out_e_bits_sink = auto_in_e_bits_sink; 
  assign TLMonitor_clock = clock; 
  assign TLMonitor_reset = reset; 
  assign TLMonitor_io_in_a_ready = _T_822 & _T_667; 
  assign TLMonitor_io_in_a_valid = auto_in_a_valid; 
  assign TLMonitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; 
  assign TLMonitor_io_in_a_bits_param = auto_in_a_bits_param; 
  assign TLMonitor_io_in_a_bits_size = auto_in_a_bits_size; 
  assign TLMonitor_io_in_a_bits_source = auto_in_a_bits_source; 
  assign TLMonitor_io_in_a_bits_address = auto_in_a_bits_address; 
  assign TLMonitor_io_in_a_bits_mask = auto_in_a_bits_mask; 
  assign TLMonitor_io_in_c_ready = auto_out_c_ready; 
  assign TLMonitor_io_in_c_valid = auto_in_c_valid; 
  assign TLMonitor_io_in_c_bits_opcode = auto_in_c_bits_opcode; 
  assign TLMonitor_io_in_c_bits_param = auto_in_c_bits_param; 
  assign TLMonitor_io_in_c_bits_size = auto_in_c_bits_size; 
  assign TLMonitor_io_in_c_bits_source = auto_in_c_bits_source; 
  assign TLMonitor_io_in_c_bits_address = auto_in_c_bits_address; 
  assign TLMonitor_io_in_c_bits_corrupt = auto_in_c_bits_corrupt; 
  assign TLMonitor_io_in_d_ready = auto_in_d_ready; 
  assign TLMonitor_io_in_d_valid = auto_out_d_valid & _T_908; 
  assign TLMonitor_io_in_d_bits_opcode = _T_907 ? 3'h1 : auto_out_d_bits_opcode; 
  assign TLMonitor_io_in_d_bits_param = auto_out_d_bits_param; 
  assign TLMonitor_io_in_d_bits_size = auto_out_d_bits_size; 
  assign TLMonitor_io_in_d_bits_source = auto_out_d_bits_source; 
  assign TLMonitor_io_in_d_bits_sink = auto_out_d_bits_sink; 
  assign TLMonitor_io_in_d_bits_denied = _T_907 ? _T_912 : auto_out_d_bits_denied; 
  assign TLMonitor_io_in_d_bits_corrupt = _T_907 ? _T_911 : auto_out_d_bits_corrupt; 
  assign TLMonitor_io_in_e_ready = auto_out_e_ready; 
  assign TLMonitor_io_in_e_valid = auto_in_e_valid; 
  assign TLMonitor_io_in_e_bits_sink = auto_in_e_bits_sink; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_10_0_state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_11_0_bits_opcode = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_11_0_bits_param = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_11_0_bits_size = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_11_0_bits_source = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_11_0_bits_address = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_11_0_bits_mask = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{`RANDOM}};
  _T_11_0_bits_data = _RAND_7[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_11_0_fifoId = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_11_0_lut = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{`RANDOM}};
  _T_12_0_data = _RAND_10[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_12_0_denied = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_12_0_corrupt = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_774 = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_818_1 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_818_0 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_883 = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_10_0_state <= 2'h0;
    end else begin
      if (_T_901) begin
        if (_T_895) begin
          if (_T_898) begin
            _T_10_0_state <= 2'h2;
          end else begin
            _T_10_0_state <= 2'h0;
          end
        end else begin
          if (_T_874) begin
            if (_T_14) begin
              _T_10_0_state <= 2'h1;
            end else begin
              if (_T_864) begin
                if (_T_13) begin
                  _T_10_0_state <= 2'h3;
                end
              end
            end
          end else begin
            if (_T_864) begin
              if (_T_13) begin
                _T_10_0_state <= 2'h3;
              end
            end
          end
        end
      end else begin
        if (_T_874) begin
          if (_T_14) begin
            _T_10_0_state <= 2'h1;
          end else begin
            if (_T_864) begin
              if (_T_13) begin
                _T_10_0_state <= 2'h3;
              end
            end
          end
        end else begin
          if (_T_864) begin
            if (_T_13) begin
              _T_10_0_state <= 2'h3;
            end
          end
        end
      end
    end
    if (_T_864) begin
      if (_T_13) begin
        _T_11_0_bits_opcode <= auto_in_a_bits_opcode;
      end
    end
    if (_T_864) begin
      if (_T_13) begin
        _T_11_0_bits_param <= auto_in_a_bits_param;
      end
    end
    if (_T_864) begin
      if (_T_13) begin
        _T_11_0_bits_size <= auto_in_a_bits_size;
      end
    end
    if (_T_864) begin
      if (_T_13) begin
        _T_11_0_bits_source <= auto_in_a_bits_source;
      end
    end
    if (_T_864) begin
      if (_T_13) begin
        _T_11_0_bits_address <= auto_in_a_bits_address;
      end
    end
    if (_T_864) begin
      if (_T_13) begin
        _T_11_0_bits_mask <= auto_in_a_bits_mask;
      end
    end
    if (_T_864) begin
      if (_T_13) begin
        _T_11_0_bits_data <= auto_in_a_bits_data;
      end
    end
    if (_T_864) begin
      if (_T_13) begin
        _T_11_0_fifoId <= _T_97;
      end
    end
    if (_T_864) begin
      if (_T_13) begin
        if (_T_872) begin
          _T_11_0_lut <= 4'h8;
        end else begin
          if (_T_870) begin
            _T_11_0_lut <= 4'he;
          end else begin
            if (_T_868) begin
              _T_11_0_lut <= 4'h6;
            end else begin
              if (_T_866) begin
                _T_11_0_lut <= 4'hc;
              end else begin
                _T_11_0_lut <= 4'h0;
              end
            end
          end
        end
      end
    end
    if (_T_901) begin
      if (_T_902) begin
        _T_12_0_data <= auto_out_d_bits_data;
      end
    end
    if (_T_901) begin
      if (_T_902) begin
        _T_12_0_denied <= auto_out_d_bits_denied;
      end
    end
    if (_T_901) begin
      if (_T_902) begin
        _T_12_0_corrupt <= auto_out_d_bits_corrupt;
      end
    end
    if (reset) begin
      _T_774 <= 5'h0;
    end else begin
      if (_T_776) begin
        if (_T_789) begin
          if (_T_772) begin
            _T_774 <= _T_770;
          end else begin
            _T_774 <= 5'h0;
          end
        end else begin
          _T_774 <= 5'h0;
        end
      end else begin
        _T_774 <= _T_815;
      end
    end
    if (reset) begin
      _T_818_1 <= 1'h0;
    end else begin
      if (_T_775) begin
        _T_818_1 <= _T_789;
      end
    end
    if (reset) begin
      _T_818_0 <= 1'h0;
    end else begin
      if (_T_775) begin
        _T_818_0 <= _T_788;
      end
    end
    if (reset) begin
      _T_883 <= 5'h0;
    end else begin
      if (_T_875) begin
        if (_T_886) begin
          if (_T_881) begin
            _T_883 <= _T_880;
          end else begin
            _T_883 <= 5'h0;
          end
        end else begin
          _T_883 <= _T_885;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_802) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_802) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_809) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:70 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_809) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLBuffer( 
  input         clock, 
  input         reset, 
  input         auto_out_c_ready, 
  output        auto_out_c_valid, 
  output [2:0]  auto_out_c_bits_opcode, 
  output [2:0]  auto_out_c_bits_param, 
  output [3:0]  auto_out_c_bits_size, 
  output        auto_out_c_bits_source, 
  output [31:0] auto_out_c_bits_address, 
  output        auto_out_c_bits_corrupt, 
  input         auto_out_d_valid, 
  input  [2:0]  auto_out_d_bits_opcode, 
  input  [1:0]  auto_out_d_bits_param, 
  input  [3:0]  auto_out_d_bits_size, 
  input         auto_out_d_bits_source, 
  input         auto_out_d_bits_sink, 
  input         auto_out_d_bits_denied, 
  input         auto_out_d_bits_corrupt 
);
  wire  TLMonitor_clock; 
  wire  TLMonitor_reset; 
  wire  TLMonitor_io_in_d_valid; 
  wire [2:0] TLMonitor_io_in_d_bits_opcode; 
  wire [1:0] TLMonitor_io_in_d_bits_param; 
  wire [3:0] TLMonitor_io_in_d_bits_size; 
  wire  TLMonitor_io_in_d_bits_source; 
  wire  TLMonitor_io_in_d_bits_sink; 
  wire  TLMonitor_io_in_d_bits_denied; 
  wire  TLMonitor_io_in_d_bits_corrupt; 
  wire  Queue_clock; 
  wire  Queue_reset; 
  wire  Queue_io_deq_ready; 
  wire  Queue_io_deq_valid; 
  wire [2:0] Queue_io_deq_bits_opcode; 
  wire [2:0] Queue_io_deq_bits_param; 
  wire [3:0] Queue_io_deq_bits_size; 
  wire  Queue_io_deq_bits_source; 
  wire [31:0] Queue_io_deq_bits_address; 
  wire  Queue_io_deq_bits_corrupt; 
  dual_TLMonitor_7 dual_TLMonitor ( 
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt)
  );
  dual_Queue_4 dual_Queue ( 
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_opcode(Queue_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_io_deq_bits_param),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_source(Queue_io_deq_bits_source),
    .io_deq_bits_address(Queue_io_deq_bits_address),
    .io_deq_bits_corrupt(Queue_io_deq_bits_corrupt)
  );
  assign auto_out_c_valid = Queue_io_deq_valid; 
  assign auto_out_c_bits_opcode = Queue_io_deq_bits_opcode; 
  assign auto_out_c_bits_param = Queue_io_deq_bits_param; 
  assign auto_out_c_bits_size = Queue_io_deq_bits_size; 
  assign auto_out_c_bits_source = Queue_io_deq_bits_source; 
  assign auto_out_c_bits_address = Queue_io_deq_bits_address; 
  assign auto_out_c_bits_corrupt = Queue_io_deq_bits_corrupt; 
  assign TLMonitor_clock = clock; 
  assign TLMonitor_reset = reset; 
  assign TLMonitor_io_in_d_valid = auto_out_d_valid; 
  assign TLMonitor_io_in_d_bits_opcode = auto_out_d_bits_opcode; 
  assign TLMonitor_io_in_d_bits_param = auto_out_d_bits_param; 
  assign TLMonitor_io_in_d_bits_size = auto_out_d_bits_size; 
  assign TLMonitor_io_in_d_bits_source = auto_out_d_bits_source; 
  assign TLMonitor_io_in_d_bits_sink = auto_out_d_bits_sink; 
  assign TLMonitor_io_in_d_bits_denied = auto_out_d_bits_denied; 
  assign TLMonitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; 
  assign Queue_clock = clock; 
  assign Queue_reset = reset; 
  assign Queue_io_deq_ready = auto_out_c_ready; 
endmodule
module dual_TLBusBypassBar( 
  input          clock, 
  input          reset, 
  output         auto_in_a_ready, 
  input          auto_in_a_valid, 
  input  [2:0]   auto_in_a_bits_opcode, 
  input  [2:0]   auto_in_a_bits_param, 
  input  [2:0]   auto_in_a_bits_size, 
  input  [2:0]   auto_in_a_bits_source, 
  input  [31:0]  auto_in_a_bits_address, 
  input  [3:0]   auto_in_a_bits_mask, 
  input  [31:0]  auto_in_a_bits_data, 
  input          auto_in_a_bits_corrupt, 
  input          auto_in_d_ready, 
  output         auto_in_d_valid, 
  output [2:0]   auto_in_d_bits_opcode, 
  output [1:0]   auto_in_d_bits_param, 
  output [2:0]   auto_in_d_bits_size, 
  output [2:0]   auto_in_d_bits_source, 
  output [4:0]   auto_in_d_bits_sink, 
  output         auto_in_d_bits_denied, 
  output [31:0]  auto_in_d_bits_data, 
  output         auto_in_d_bits_corrupt, 
  input          auto_out_1_a_ready, 
  output         auto_out_1_a_valid, 
  output [2:0]   auto_out_1_a_bits_opcode, 
  output [2:0]   auto_out_1_a_bits_param, 
  output [2:0]   auto_out_1_a_bits_size, 
  output [2:0]   auto_out_1_a_bits_source, 
  output [31:0]  auto_out_1_a_bits_address, 
  output [3:0]   auto_out_1_a_bits_mask, 
  output [31:0]  auto_out_1_a_bits_data, 
  output         auto_out_1_a_bits_corrupt, 
  output         auto_out_1_d_ready, 
  input          auto_out_1_d_valid, 
  input  [2:0]   auto_out_1_d_bits_opcode, 
  input  [1:0]   auto_out_1_d_bits_param, 
  input  [2:0]   auto_out_1_d_bits_size, 
  input  [2:0]   auto_out_1_d_bits_source, 
  input  [4:0]   auto_out_1_d_bits_sink, 
  input          auto_out_1_d_bits_denied, 
  input  [31:0]  auto_out_1_d_bits_data, 
  input          auto_out_1_d_bits_corrupt, 
  input          auto_out_0_a_ready, 
  output         auto_out_0_a_valid, 
  output [2:0]   auto_out_0_a_bits_opcode, 
  output [2:0]   auto_out_0_a_bits_param, 
  output [3:0]   auto_out_0_a_bits_size, 
  output [2:0]   auto_out_0_a_bits_source, 
  output [127:0] auto_out_0_a_bits_address, 
  output [3:0]   auto_out_0_a_bits_mask, 
  output         auto_out_0_a_bits_corrupt, 
  output         auto_out_0_d_ready, 
  input          auto_out_0_d_valid, 
  input  [2:0]   auto_out_0_d_bits_opcode, 
  input  [1:0]   auto_out_0_d_bits_param, 
  input  [3:0]   auto_out_0_d_bits_size, 
  input  [2:0]   auto_out_0_d_bits_source, 
  input          auto_out_0_d_bits_sink, 
  input          auto_out_0_d_bits_denied, 
  input  [31:0]  auto_out_0_d_bits_data, 
  input          auto_out_0_d_bits_corrupt, 
  input          io_bypass 
);
  wire  TLMonitor_clock; 
  wire  TLMonitor_reset; 
  wire  TLMonitor_io_in_a_ready; 
  wire  TLMonitor_io_in_a_valid; 
  wire [2:0] TLMonitor_io_in_a_bits_opcode; 
  wire [2:0] TLMonitor_io_in_a_bits_param; 
  wire [2:0] TLMonitor_io_in_a_bits_size; 
  wire [2:0] TLMonitor_io_in_a_bits_source; 
  wire [31:0] TLMonitor_io_in_a_bits_address; 
  wire [3:0] TLMonitor_io_in_a_bits_mask; 
  wire  TLMonitor_io_in_a_bits_corrupt; 
  wire  TLMonitor_io_in_d_ready; 
  wire  TLMonitor_io_in_d_valid; 
  wire [2:0] TLMonitor_io_in_d_bits_opcode; 
  wire [1:0] TLMonitor_io_in_d_bits_param; 
  wire [2:0] TLMonitor_io_in_d_bits_size; 
  wire [2:0] TLMonitor_io_in_d_bits_source; 
  wire [4:0] TLMonitor_io_in_d_bits_sink; 
  wire  TLMonitor_io_in_d_bits_denied; 
  wire  TLMonitor_io_in_d_bits_corrupt; 
  reg  bypass; 
  reg [31:0] _RAND_0;
  reg [4:0] flight; 
  reg [31:0] _RAND_1;
  wire  _T_151; 
  reg [3:0] _T_161; 
  reg [31:0] _RAND_2;
  wire  _T_164; 
  wire  stall; 
  wire  _T_179; 
  wire  _T_180; 
  wire  in_a_ready; 
  wire  _T_6; 
  wire [12:0] _T_8; 
  wire [5:0] _T_9; 
  wire [5:0] _T_10; 
  wire [3:0] _T_11; 
  wire  _T_12; 
  wire  _T_13; 
  reg [3:0] _T_15; 
  reg [31:0] _RAND_3;
  wire [3:0] _T_17; 
  wire  _T_18; 
  wire  in_d_valid; 
  wire  _T_65; 
  wire [2:0] _T_186_size; 
  wire [2:0] in_d_bits_size; 
  wire [12:0] _T_67; 
  wire [5:0] _T_68; 
  wire [5:0] _T_69; 
  wire [3:0] _T_70; 
  wire [2:0] in_d_bits_opcode; 
  wire  _T_71; 
  wire [3:0] _T_72; 
  reg [3:0] _T_73; 
  reg [31:0] _RAND_4;
  wire [3:0] _T_75; 
  wire  _T_76; 
  wire  _T_77; 
  wire  _T_78; 
  wire  _T_79; 
  wire  _T_104; 
  wire  _T_105; 
  wire  _T_106; 
  wire  _T_107; 
  wire  _T_109; 
  wire  _T_118; 
  wire  _T_119; 
  wire [1:0] _T_123; 
  wire  _T_134; 
  wire [1:0] _T_139; 
  wire  _T_140; 
  wire  _T_141; 
  wire [1:0] _T_142; 
  wire [4:0] _GEN_7; 
  wire [4:0] _T_144; 
  wire  _T_145; 
  wire  _T_146; 
  wire [1:0] _T_147; 
  wire [4:0] _GEN_8; 
  wire [4:0] next_flight; 
  wire  _T_150; 
  wire [3:0] _T_163; 
  wire  _T_173; 
  wire  _T_177; 
  wire [4:0] _T_186_sink; 
  dual_TLMonitor_3 dual_TLMonitor ( 
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_io_in_a_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt)
  );
  assign _T_151 = bypass != io_bypass; 
  assign _T_164 = _T_161 == 4'h0; 
  assign stall = _T_151 & _T_164; 
  assign _T_179 = stall == 1'h0; 
  assign _T_180 = bypass ? auto_out_0_a_ready : auto_out_1_a_ready; 
  assign in_a_ready = _T_179 & _T_180; 
  assign _T_6 = in_a_ready & auto_in_a_valid; 
  assign _T_8 = 13'h3f << auto_in_a_bits_size; 
  assign _T_9 = _T_8[5:0]; 
  assign _T_10 = ~ _T_9; 
  assign _T_11 = _T_10[5:2]; 
  assign _T_12 = auto_in_a_bits_opcode[2]; 
  assign _T_13 = _T_12 == 1'h0; 
  assign _T_17 = _T_15 - 4'h1; 
  assign _T_18 = _T_15 == 4'h0; 
  assign in_d_valid = bypass ? auto_out_0_d_valid : auto_out_1_d_valid; 
  assign _T_65 = auto_in_d_ready & in_d_valid; 
  assign _T_186_size = auto_out_0_d_bits_size[2:0]; 
  assign in_d_bits_size = bypass ? _T_186_size : auto_out_1_d_bits_size; 
  assign _T_67 = 13'h3f << in_d_bits_size; 
  assign _T_68 = _T_67[5:0]; 
  assign _T_69 = ~ _T_68; 
  assign _T_70 = _T_69[5:2]; 
  assign in_d_bits_opcode = bypass ? auto_out_0_d_bits_opcode : auto_out_1_d_bits_opcode; 
  assign _T_71 = in_d_bits_opcode[0]; 
  assign _T_72 = _T_71 ? _T_70 : 4'h0; 
  assign _T_75 = _T_73 - 4'h1; 
  assign _T_76 = _T_73 == 4'h0; 
  assign _T_77 = _T_73 == 4'h1; 
  assign _T_78 = _T_72 == 4'h0; 
  assign _T_79 = _T_77 | _T_78; 
  assign _T_104 = in_d_bits_opcode[2]; 
  assign _T_105 = in_d_bits_opcode[1]; 
  assign _T_106 = _T_105 == 1'h0; 
  assign _T_107 = _T_104 & _T_106; 
  assign _T_109 = _T_6 & _T_18; 
  assign _T_118 = _T_65 & _T_76; 
  assign _T_119 = _T_118 & _T_107; 
  assign _T_123 = {_T_109,_T_119}; 
  assign _T_134 = _T_65 & _T_79; 
  assign _T_139 = {1'h0,_T_134}; 
  assign _T_140 = _T_123[0]; 
  assign _T_141 = _T_123[1]; 
  assign _T_142 = _T_140 + _T_141; 
  assign _GEN_7 = {{3'd0}, _T_142}; 
  assign _T_144 = flight + _GEN_7; 
  assign _T_145 = _T_139[0]; 
  assign _T_146 = _T_139[1]; 
  assign _T_147 = _T_145 + _T_146; 
  assign _GEN_8 = {{3'd0}, _T_147}; 
  assign next_flight = _T_144 - _GEN_8; 
  assign _T_150 = next_flight == 5'h0; 
  assign _T_163 = _T_161 - 4'h1; 
  assign _T_173 = _T_179 & auto_in_a_valid; 
  assign _T_177 = bypass == 1'h0; 
  assign _T_186_sink = {{4'd0}, auto_out_0_d_bits_sink}; 
  assign auto_in_a_ready = _T_179 & _T_180; 
  assign auto_in_d_valid = bypass ? auto_out_0_d_valid : auto_out_1_d_valid; 
  assign auto_in_d_bits_opcode = bypass ? auto_out_0_d_bits_opcode : auto_out_1_d_bits_opcode; 
  assign auto_in_d_bits_param = bypass ? auto_out_0_d_bits_param : auto_out_1_d_bits_param; 
  assign auto_in_d_bits_size = bypass ? _T_186_size : auto_out_1_d_bits_size; 
  assign auto_in_d_bits_source = bypass ? auto_out_0_d_bits_source : auto_out_1_d_bits_source; 
  assign auto_in_d_bits_sink = bypass ? _T_186_sink : auto_out_1_d_bits_sink; 
  assign auto_in_d_bits_denied = bypass ? auto_out_0_d_bits_denied : auto_out_1_d_bits_denied; 
  assign auto_in_d_bits_data = bypass ? auto_out_0_d_bits_data : auto_out_1_d_bits_data; 
  assign auto_in_d_bits_corrupt = bypass ? auto_out_0_d_bits_corrupt : auto_out_1_d_bits_corrupt; 
  assign auto_out_1_a_valid = _T_173 & _T_177; 
  assign auto_out_1_a_bits_opcode = auto_in_a_bits_opcode; 
  assign auto_out_1_a_bits_param = auto_in_a_bits_param; 
  assign auto_out_1_a_bits_size = auto_in_a_bits_size; 
  assign auto_out_1_a_bits_source = auto_in_a_bits_source; 
  assign auto_out_1_a_bits_address = auto_in_a_bits_address; 
  assign auto_out_1_a_bits_mask = auto_in_a_bits_mask; 
  assign auto_out_1_a_bits_data = auto_in_a_bits_data; 
  assign auto_out_1_a_bits_corrupt = auto_in_a_bits_corrupt; 
  assign auto_out_1_d_ready = auto_in_d_ready & _T_177; 
  assign auto_out_0_a_valid = _T_173 & bypass; 
  assign auto_out_0_a_bits_opcode = auto_in_a_bits_opcode; 
  assign auto_out_0_a_bits_param = auto_in_a_bits_param; 
  assign auto_out_0_a_bits_size = {{1'd0}, auto_in_a_bits_size}; 
  assign auto_out_0_a_bits_source = auto_in_a_bits_source; 
  assign auto_out_0_a_bits_address = {{96'd0}, auto_in_a_bits_address}; 
  assign auto_out_0_a_bits_mask = auto_in_a_bits_mask; 
  assign auto_out_0_a_bits_corrupt = auto_in_a_bits_corrupt; 
  assign auto_out_0_d_ready = auto_in_d_ready & bypass; 
  assign TLMonitor_clock = clock; 
  assign TLMonitor_reset = reset; 
  assign TLMonitor_io_in_a_ready = _T_179 & _T_180; 
  assign TLMonitor_io_in_a_valid = auto_in_a_valid; 
  assign TLMonitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; 
  assign TLMonitor_io_in_a_bits_param = auto_in_a_bits_param; 
  assign TLMonitor_io_in_a_bits_size = auto_in_a_bits_size; 
  assign TLMonitor_io_in_a_bits_source = auto_in_a_bits_source; 
  assign TLMonitor_io_in_a_bits_address = auto_in_a_bits_address; 
  assign TLMonitor_io_in_a_bits_mask = auto_in_a_bits_mask; 
  assign TLMonitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; 
  assign TLMonitor_io_in_d_ready = auto_in_d_ready; 
  assign TLMonitor_io_in_d_valid = bypass ? auto_out_0_d_valid : auto_out_1_d_valid; 
  assign TLMonitor_io_in_d_bits_opcode = bypass ? auto_out_0_d_bits_opcode : auto_out_1_d_bits_opcode; 
  assign TLMonitor_io_in_d_bits_param = bypass ? auto_out_0_d_bits_param : auto_out_1_d_bits_param; 
  assign TLMonitor_io_in_d_bits_size = bypass ? _T_186_size : auto_out_1_d_bits_size; 
  assign TLMonitor_io_in_d_bits_source = bypass ? auto_out_0_d_bits_source : auto_out_1_d_bits_source; 
  assign TLMonitor_io_in_d_bits_sink = bypass ? _T_186_sink : auto_out_1_d_bits_sink; 
  assign TLMonitor_io_in_d_bits_denied = bypass ? auto_out_0_d_bits_denied : auto_out_1_d_bits_denied; 
  assign TLMonitor_io_in_d_bits_corrupt = bypass ? auto_out_0_d_bits_corrupt : auto_out_1_d_bits_corrupt; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bypass = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  flight = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_161 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_15 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_73 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      bypass <= io_bypass;
    end else begin
      if (_T_150) begin
        bypass <= io_bypass;
      end
    end
    if (reset) begin
      flight <= 5'h0;
    end else begin
      flight <= next_flight;
    end
    if (reset) begin
      _T_161 <= 4'h0;
    end else begin
      if (_T_6) begin
        if (_T_164) begin
          if (_T_13) begin
            _T_161 <= _T_11;
          end else begin
            _T_161 <= 4'h0;
          end
        end else begin
          _T_161 <= _T_163;
        end
      end
    end
    if (reset) begin
      _T_15 <= 4'h0;
    end else begin
      if (_T_6) begin
        if (_T_18) begin
          if (_T_13) begin
            _T_15 <= _T_11;
          end else begin
            _T_15 <= 4'h0;
          end
        end else begin
          _T_15 <= _T_17;
        end
      end
    end
    if (reset) begin
      _T_73 <= 4'h0;
    end else begin
      if (_T_65) begin
        if (_T_76) begin
          if (_T_71) begin
            _T_73 <= _T_70;
          end else begin
            _T_73 <= 4'h0;
          end
        end else begin
          _T_73 <= _T_75;
        end
      end
    end
  end
endmodule
module dual_TLBusBypass( 
  input         clock, 
  input         reset, 
  input         auto_node_out_out_a_ready, 
  output        auto_node_out_out_a_valid, 
  output [2:0]  auto_node_out_out_a_bits_opcode, 
  output [2:0]  auto_node_out_out_a_bits_param, 
  output [2:0]  auto_node_out_out_a_bits_size, 
  output [2:0]  auto_node_out_out_a_bits_source, 
  output [31:0] auto_node_out_out_a_bits_address, 
  output [3:0]  auto_node_out_out_a_bits_mask, 
  output [31:0] auto_node_out_out_a_bits_data, 
  output        auto_node_out_out_a_bits_corrupt, 
  output        auto_node_out_out_d_ready, 
  input         auto_node_out_out_d_valid, 
  input  [2:0]  auto_node_out_out_d_bits_opcode, 
  input  [1:0]  auto_node_out_out_d_bits_param, 
  input  [2:0]  auto_node_out_out_d_bits_size, 
  input  [2:0]  auto_node_out_out_d_bits_source, 
  input  [4:0]  auto_node_out_out_d_bits_sink, 
  input         auto_node_out_out_d_bits_denied, 
  input  [31:0] auto_node_out_out_d_bits_data, 
  input         auto_node_out_out_d_bits_corrupt, 
  output        auto_node_in_in_a_ready, 
  input         auto_node_in_in_a_valid, 
  input  [2:0]  auto_node_in_in_a_bits_opcode, 
  input  [2:0]  auto_node_in_in_a_bits_param, 
  input  [2:0]  auto_node_in_in_a_bits_size, 
  input  [2:0]  auto_node_in_in_a_bits_source, 
  input  [31:0] auto_node_in_in_a_bits_address, 
  input  [3:0]  auto_node_in_in_a_bits_mask, 
  input  [31:0] auto_node_in_in_a_bits_data, 
  input         auto_node_in_in_a_bits_corrupt, 
  input         auto_node_in_in_d_ready, 
  output        auto_node_in_in_d_valid, 
  output [2:0]  auto_node_in_in_d_bits_opcode, 
  output [1:0]  auto_node_in_in_d_bits_param, 
  output [2:0]  auto_node_in_in_d_bits_size, 
  output [2:0]  auto_node_in_in_d_bits_source, 
  output [4:0]  auto_node_in_in_d_bits_sink, 
  output        auto_node_in_in_d_bits_denied, 
  output [31:0] auto_node_in_in_d_bits_data, 
  output        auto_node_in_in_d_bits_corrupt, 
  input         io_bypass 
);
  wire  bar_clock; 
  wire  bar_reset; 
  wire  bar_auto_in_a_ready; 
  wire  bar_auto_in_a_valid; 
  wire [2:0] bar_auto_in_a_bits_opcode; 
  wire [2:0] bar_auto_in_a_bits_param; 
  wire [2:0] bar_auto_in_a_bits_size; 
  wire [2:0] bar_auto_in_a_bits_source; 
  wire [31:0] bar_auto_in_a_bits_address; 
  wire [3:0] bar_auto_in_a_bits_mask; 
  wire [31:0] bar_auto_in_a_bits_data; 
  wire  bar_auto_in_a_bits_corrupt; 
  wire  bar_auto_in_d_ready; 
  wire  bar_auto_in_d_valid; 
  wire [2:0] bar_auto_in_d_bits_opcode; 
  wire [1:0] bar_auto_in_d_bits_param; 
  wire [2:0] bar_auto_in_d_bits_size; 
  wire [2:0] bar_auto_in_d_bits_source; 
  wire [4:0] bar_auto_in_d_bits_sink; 
  wire  bar_auto_in_d_bits_denied; 
  wire [31:0] bar_auto_in_d_bits_data; 
  wire  bar_auto_in_d_bits_corrupt; 
  wire  bar_auto_out_1_a_ready; 
  wire  bar_auto_out_1_a_valid; 
  wire [2:0] bar_auto_out_1_a_bits_opcode; 
  wire [2:0] bar_auto_out_1_a_bits_param; 
  wire [2:0] bar_auto_out_1_a_bits_size; 
  wire [2:0] bar_auto_out_1_a_bits_source; 
  wire [31:0] bar_auto_out_1_a_bits_address; 
  wire [3:0] bar_auto_out_1_a_bits_mask; 
  wire [31:0] bar_auto_out_1_a_bits_data; 
  wire  bar_auto_out_1_a_bits_corrupt; 
  wire  bar_auto_out_1_d_ready; 
  wire  bar_auto_out_1_d_valid; 
  wire [2:0] bar_auto_out_1_d_bits_opcode; 
  wire [1:0] bar_auto_out_1_d_bits_param; 
  wire [2:0] bar_auto_out_1_d_bits_size; 
  wire [2:0] bar_auto_out_1_d_bits_source; 
  wire [4:0] bar_auto_out_1_d_bits_sink; 
  wire  bar_auto_out_1_d_bits_denied; 
  wire [31:0] bar_auto_out_1_d_bits_data; 
  wire  bar_auto_out_1_d_bits_corrupt; 
  wire  bar_auto_out_0_a_ready; 
  wire  bar_auto_out_0_a_valid; 
  wire [2:0] bar_auto_out_0_a_bits_opcode; 
  wire [2:0] bar_auto_out_0_a_bits_param; 
  wire [3:0] bar_auto_out_0_a_bits_size; 
  wire [2:0] bar_auto_out_0_a_bits_source; 
  wire [127:0] bar_auto_out_0_a_bits_address; 
  wire [3:0] bar_auto_out_0_a_bits_mask; 
  wire  bar_auto_out_0_a_bits_corrupt; 
  wire  bar_auto_out_0_d_ready; 
  wire  bar_auto_out_0_d_valid; 
  wire [2:0] bar_auto_out_0_d_bits_opcode; 
  wire [1:0] bar_auto_out_0_d_bits_param; 
  wire [3:0] bar_auto_out_0_d_bits_size; 
  wire [2:0] bar_auto_out_0_d_bits_source; 
  wire  bar_auto_out_0_d_bits_sink; 
  wire  bar_auto_out_0_d_bits_denied; 
  wire [31:0] bar_auto_out_0_d_bits_data; 
  wire  bar_auto_out_0_d_bits_corrupt; 
  wire  bar_io_bypass; 
  wire  error_clock; 
  wire  error_reset; 
  wire  error_auto_in_a_ready; 
  wire  error_auto_in_a_valid; 
  wire [2:0] error_auto_in_a_bits_opcode; 
  wire [2:0] error_auto_in_a_bits_param; 
  wire [3:0] error_auto_in_a_bits_size; 
  wire [2:0] error_auto_in_a_bits_source; 
  wire [127:0] error_auto_in_a_bits_address; 
  wire [3:0] error_auto_in_a_bits_mask; 
  wire  error_auto_in_a_bits_corrupt; 
  wire  error_auto_in_d_ready; 
  wire  error_auto_in_d_valid; 
  wire [2:0] error_auto_in_d_bits_opcode; 
  wire [1:0] error_auto_in_d_bits_param; 
  wire [3:0] error_auto_in_d_bits_size; 
  wire [2:0] error_auto_in_d_bits_source; 
  wire  error_auto_in_d_bits_sink; 
  wire  error_auto_in_d_bits_denied; 
  wire [31:0] error_auto_in_d_bits_data; 
  wire  error_auto_in_d_bits_corrupt; 
  dual_TLBusBypassBar bar ( 
    .clock(bar_clock),
    .reset(bar_reset),
    .auto_in_a_ready(bar_auto_in_a_ready),
    .auto_in_a_valid(bar_auto_in_a_valid),
    .auto_in_a_bits_opcode(bar_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(bar_auto_in_a_bits_param),
    .auto_in_a_bits_size(bar_auto_in_a_bits_size),
    .auto_in_a_bits_source(bar_auto_in_a_bits_source),
    .auto_in_a_bits_address(bar_auto_in_a_bits_address),
    .auto_in_a_bits_mask(bar_auto_in_a_bits_mask),
    .auto_in_a_bits_data(bar_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(bar_auto_in_a_bits_corrupt),
    .auto_in_d_ready(bar_auto_in_d_ready),
    .auto_in_d_valid(bar_auto_in_d_valid),
    .auto_in_d_bits_opcode(bar_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(bar_auto_in_d_bits_param),
    .auto_in_d_bits_size(bar_auto_in_d_bits_size),
    .auto_in_d_bits_source(bar_auto_in_d_bits_source),
    .auto_in_d_bits_sink(bar_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(bar_auto_in_d_bits_denied),
    .auto_in_d_bits_data(bar_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(bar_auto_in_d_bits_corrupt),
    .auto_out_1_a_ready(bar_auto_out_1_a_ready),
    .auto_out_1_a_valid(bar_auto_out_1_a_valid),
    .auto_out_1_a_bits_opcode(bar_auto_out_1_a_bits_opcode),
    .auto_out_1_a_bits_param(bar_auto_out_1_a_bits_param),
    .auto_out_1_a_bits_size(bar_auto_out_1_a_bits_size),
    .auto_out_1_a_bits_source(bar_auto_out_1_a_bits_source),
    .auto_out_1_a_bits_address(bar_auto_out_1_a_bits_address),
    .auto_out_1_a_bits_mask(bar_auto_out_1_a_bits_mask),
    .auto_out_1_a_bits_data(bar_auto_out_1_a_bits_data),
    .auto_out_1_a_bits_corrupt(bar_auto_out_1_a_bits_corrupt),
    .auto_out_1_d_ready(bar_auto_out_1_d_ready),
    .auto_out_1_d_valid(bar_auto_out_1_d_valid),
    .auto_out_1_d_bits_opcode(bar_auto_out_1_d_bits_opcode),
    .auto_out_1_d_bits_param(bar_auto_out_1_d_bits_param),
    .auto_out_1_d_bits_size(bar_auto_out_1_d_bits_size),
    .auto_out_1_d_bits_source(bar_auto_out_1_d_bits_source),
    .auto_out_1_d_bits_sink(bar_auto_out_1_d_bits_sink),
    .auto_out_1_d_bits_denied(bar_auto_out_1_d_bits_denied),
    .auto_out_1_d_bits_data(bar_auto_out_1_d_bits_data),
    .auto_out_1_d_bits_corrupt(bar_auto_out_1_d_bits_corrupt),
    .auto_out_0_a_ready(bar_auto_out_0_a_ready),
    .auto_out_0_a_valid(bar_auto_out_0_a_valid),
    .auto_out_0_a_bits_opcode(bar_auto_out_0_a_bits_opcode),
    .auto_out_0_a_bits_param(bar_auto_out_0_a_bits_param),
    .auto_out_0_a_bits_size(bar_auto_out_0_a_bits_size),
    .auto_out_0_a_bits_source(bar_auto_out_0_a_bits_source),
    .auto_out_0_a_bits_address(bar_auto_out_0_a_bits_address),
    .auto_out_0_a_bits_mask(bar_auto_out_0_a_bits_mask),
    .auto_out_0_a_bits_corrupt(bar_auto_out_0_a_bits_corrupt),
    .auto_out_0_d_ready(bar_auto_out_0_d_ready),
    .auto_out_0_d_valid(bar_auto_out_0_d_valid),
    .auto_out_0_d_bits_opcode(bar_auto_out_0_d_bits_opcode),
    .auto_out_0_d_bits_param(bar_auto_out_0_d_bits_param),
    .auto_out_0_d_bits_size(bar_auto_out_0_d_bits_size),
    .auto_out_0_d_bits_source(bar_auto_out_0_d_bits_source),
    .auto_out_0_d_bits_sink(bar_auto_out_0_d_bits_sink),
    .auto_out_0_d_bits_denied(bar_auto_out_0_d_bits_denied),
    .auto_out_0_d_bits_data(bar_auto_out_0_d_bits_data),
    .auto_out_0_d_bits_corrupt(bar_auto_out_0_d_bits_corrupt),
    .io_bypass(bar_io_bypass)
  );
  dual_TLError_1 error ( 
    .clock(error_clock),
    .reset(error_reset),
    .auto_in_a_ready(error_auto_in_a_ready),
    .auto_in_a_valid(error_auto_in_a_valid),
    .auto_in_a_bits_opcode(error_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(error_auto_in_a_bits_param),
    .auto_in_a_bits_size(error_auto_in_a_bits_size),
    .auto_in_a_bits_source(error_auto_in_a_bits_source),
    .auto_in_a_bits_address(error_auto_in_a_bits_address),
    .auto_in_a_bits_mask(error_auto_in_a_bits_mask),
    .auto_in_a_bits_corrupt(error_auto_in_a_bits_corrupt),
    .auto_in_d_ready(error_auto_in_d_ready),
    .auto_in_d_valid(error_auto_in_d_valid),
    .auto_in_d_bits_opcode(error_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(error_auto_in_d_bits_param),
    .auto_in_d_bits_size(error_auto_in_d_bits_size),
    .auto_in_d_bits_source(error_auto_in_d_bits_source),
    .auto_in_d_bits_sink(error_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(error_auto_in_d_bits_denied),
    .auto_in_d_bits_data(error_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(error_auto_in_d_bits_corrupt)
  );
  assign auto_node_out_out_a_valid = bar_auto_out_1_a_valid; 
  assign auto_node_out_out_a_bits_opcode = bar_auto_out_1_a_bits_opcode; 
  assign auto_node_out_out_a_bits_param = bar_auto_out_1_a_bits_param; 
  assign auto_node_out_out_a_bits_size = bar_auto_out_1_a_bits_size; 
  assign auto_node_out_out_a_bits_source = bar_auto_out_1_a_bits_source; 
  assign auto_node_out_out_a_bits_address = bar_auto_out_1_a_bits_address; 
  assign auto_node_out_out_a_bits_mask = bar_auto_out_1_a_bits_mask; 
  assign auto_node_out_out_a_bits_data = bar_auto_out_1_a_bits_data; 
  assign auto_node_out_out_a_bits_corrupt = bar_auto_out_1_a_bits_corrupt; 
  assign auto_node_out_out_d_ready = bar_auto_out_1_d_ready; 
  assign auto_node_in_in_a_ready = bar_auto_in_a_ready; 
  assign auto_node_in_in_d_valid = bar_auto_in_d_valid; 
  assign auto_node_in_in_d_bits_opcode = bar_auto_in_d_bits_opcode; 
  assign auto_node_in_in_d_bits_param = bar_auto_in_d_bits_param; 
  assign auto_node_in_in_d_bits_size = bar_auto_in_d_bits_size; 
  assign auto_node_in_in_d_bits_source = bar_auto_in_d_bits_source; 
  assign auto_node_in_in_d_bits_sink = bar_auto_in_d_bits_sink; 
  assign auto_node_in_in_d_bits_denied = bar_auto_in_d_bits_denied; 
  assign auto_node_in_in_d_bits_data = bar_auto_in_d_bits_data; 
  assign auto_node_in_in_d_bits_corrupt = bar_auto_in_d_bits_corrupt; 
  assign bar_clock = clock; 
  assign bar_reset = reset; 
  assign bar_auto_in_a_valid = auto_node_in_in_a_valid; 
  assign bar_auto_in_a_bits_opcode = auto_node_in_in_a_bits_opcode; 
  assign bar_auto_in_a_bits_param = auto_node_in_in_a_bits_param; 
  assign bar_auto_in_a_bits_size = auto_node_in_in_a_bits_size; 
  assign bar_auto_in_a_bits_source = auto_node_in_in_a_bits_source; 
  assign bar_auto_in_a_bits_address = auto_node_in_in_a_bits_address; 
  assign bar_auto_in_a_bits_mask = auto_node_in_in_a_bits_mask; 
  assign bar_auto_in_a_bits_data = auto_node_in_in_a_bits_data; 
  assign bar_auto_in_a_bits_corrupt = auto_node_in_in_a_bits_corrupt; 
  assign bar_auto_in_d_ready = auto_node_in_in_d_ready; 
  assign bar_auto_out_1_a_ready = auto_node_out_out_a_ready; 
  assign bar_auto_out_1_d_valid = auto_node_out_out_d_valid; 
  assign bar_auto_out_1_d_bits_opcode = auto_node_out_out_d_bits_opcode; 
  assign bar_auto_out_1_d_bits_param = auto_node_out_out_d_bits_param; 
  assign bar_auto_out_1_d_bits_size = auto_node_out_out_d_bits_size; 
  assign bar_auto_out_1_d_bits_source = auto_node_out_out_d_bits_source; 
  assign bar_auto_out_1_d_bits_sink = auto_node_out_out_d_bits_sink; 
  assign bar_auto_out_1_d_bits_denied = auto_node_out_out_d_bits_denied; 
  assign bar_auto_out_1_d_bits_data = auto_node_out_out_d_bits_data; 
  assign bar_auto_out_1_d_bits_corrupt = auto_node_out_out_d_bits_corrupt; 
  assign bar_auto_out_0_a_ready = error_auto_in_a_ready; 
  assign bar_auto_out_0_d_valid = error_auto_in_d_valid; 
  assign bar_auto_out_0_d_bits_opcode = error_auto_in_d_bits_opcode; 
  assign bar_auto_out_0_d_bits_param = error_auto_in_d_bits_param; 
  assign bar_auto_out_0_d_bits_size = error_auto_in_d_bits_size; 
  assign bar_auto_out_0_d_bits_source = error_auto_in_d_bits_source; 
  assign bar_auto_out_0_d_bits_sink = error_auto_in_d_bits_sink; 
  assign bar_auto_out_0_d_bits_denied = error_auto_in_d_bits_denied; 
  assign bar_auto_out_0_d_bits_data = error_auto_in_d_bits_data; 
  assign bar_auto_out_0_d_bits_corrupt = error_auto_in_d_bits_corrupt; 
  assign bar_io_bypass = io_bypass; 
  assign error_clock = clock; 
  assign error_reset = reset; 
  assign error_auto_in_a_valid = bar_auto_out_0_a_valid; 
  assign error_auto_in_a_bits_opcode = bar_auto_out_0_a_bits_opcode; 
  assign error_auto_in_a_bits_param = bar_auto_out_0_a_bits_param; 
  assign error_auto_in_a_bits_size = bar_auto_out_0_a_bits_size; 
  assign error_auto_in_a_bits_source = bar_auto_out_0_a_bits_source; 
  assign error_auto_in_a_bits_address = bar_auto_out_0_a_bits_address; 
  assign error_auto_in_a_bits_mask = bar_auto_out_0_a_bits_mask; 
  assign error_auto_in_a_bits_corrupt = bar_auto_out_0_a_bits_corrupt; 
  assign error_auto_in_d_ready = bar_auto_out_0_d_ready; 
endmodule
module dual_TLError_1( 
  input          clock, 
  input          reset, 
  output         auto_in_a_ready, 
  input          auto_in_a_valid, 
  input  [2:0]   auto_in_a_bits_opcode, 
  input  [2:0]   auto_in_a_bits_param, 
  input  [3:0]   auto_in_a_bits_size, 
  input  [2:0]   auto_in_a_bits_source, 
  input  [127:0] auto_in_a_bits_address, 
  input  [3:0]   auto_in_a_bits_mask, 
  input          auto_in_a_bits_corrupt, 
  input          auto_in_d_ready, 
  output         auto_in_d_valid, 
  output [2:0]   auto_in_d_bits_opcode, 
  output [1:0]   auto_in_d_bits_param, 
  output [3:0]   auto_in_d_bits_size, 
  output [2:0]   auto_in_d_bits_source, 
  output         auto_in_d_bits_sink, 
  output         auto_in_d_bits_denied, 
  output [31:0]  auto_in_d_bits_data, 
  output         auto_in_d_bits_corrupt 
);
  wire  TLMonitor_clock; 
  wire  TLMonitor_reset; 
  wire  TLMonitor_io_in_a_ready; 
  wire  TLMonitor_io_in_a_valid; 
  wire [2:0] TLMonitor_io_in_a_bits_opcode; 
  wire [2:0] TLMonitor_io_in_a_bits_param; 
  wire [3:0] TLMonitor_io_in_a_bits_size; 
  wire [2:0] TLMonitor_io_in_a_bits_source; 
  wire [127:0] TLMonitor_io_in_a_bits_address; 
  wire [3:0] TLMonitor_io_in_a_bits_mask; 
  wire  TLMonitor_io_in_a_bits_corrupt; 
  wire  TLMonitor_io_in_d_ready; 
  wire  TLMonitor_io_in_d_valid; 
  wire [2:0] TLMonitor_io_in_d_bits_opcode; 
  wire [1:0] TLMonitor_io_in_d_bits_param; 
  wire [3:0] TLMonitor_io_in_d_bits_size; 
  wire [2:0] TLMonitor_io_in_d_bits_source; 
  wire  TLMonitor_io_in_d_bits_sink; 
  wire  TLMonitor_io_in_d_bits_denied; 
  wire  TLMonitor_io_in_d_bits_corrupt; 
  wire  a_clock; 
  wire  a_reset; 
  wire  a_io_enq_ready; 
  wire  a_io_enq_valid; 
  wire [2:0] a_io_enq_bits_opcode; 
  wire [3:0] a_io_enq_bits_size; 
  wire [2:0] a_io_enq_bits_source; 
  wire  a_io_deq_ready; 
  wire  a_io_deq_valid; 
  wire [2:0] a_io_deq_bits_opcode; 
  wire [3:0] a_io_deq_bits_size; 
  wire [2:0] a_io_deq_bits_source; 
  reg  idle; 
  reg [31:0] _RAND_0;
  wire  _T_6; 
  wire [26:0] _T_8; 
  wire [11:0] _T_9; 
  wire [11:0] _T_10; 
  wire [9:0] _T_11; 
  wire  _T_12; 
  wire  _T_13; 
  wire [9:0] _T_14; 
  reg [9:0] _T_15; 
  reg [31:0] _RAND_1;
  wire [9:0] _T_17; 
  wire  _T_18; 
  wire  _T_19; 
  wire  _T_20; 
  wire  a_last; 
  reg [9:0] _T_117; 
  reg [31:0] _RAND_2;
  wire  _T_118; 
  wire  _T_50; 
  wire  da_valid; 
  wire [1:0] _T_120; 
  wire [2:0] _T_121; 
  wire [1:0] _T_122; 
  wire [1:0] _T_123; 
  wire [2:0] _T_125; 
  wire [1:0] _T_126; 
  wire [1:0] _T_127; 
  wire  _T_129; 
  reg  _T_161_1; 
  reg [31:0] _RAND_3;
  wire  _T_163_1; 
  wire  da_ready; 
  wire  _T_25; 
  wire [3:0] da_bits_size; 
  wire [26:0] _T_27; 
  wire [11:0] _T_28; 
  wire [11:0] _T_29; 
  wire [9:0] _T_30; 
  wire [2:0] _GEN_4; 
  wire [2:0] _GEN_5; 
  wire [2:0] _GEN_6; 
  wire [2:0] _GEN_7; 
  wire [2:0] _GEN_8; 
  wire [2:0] da_bits_opcode; 
  wire  _T_31; 
  wire [9:0] _T_32; 
  reg [9:0] _T_33; 
  reg [31:0] _RAND_4;
  wire [9:0] _T_35; 
  wire  da_first; 
  wire  _T_36; 
  wire  _T_37; 
  wire  da_last; 
  wire  _T_42; 
  wire  _T_44; 
  wire  _T_45; 
  wire  _T_46; 
  wire  _T_47; 
  wire  _T_48; 
  wire  _T_94; 
  wire  _T_95; 
  wire  _T_119; 
  wire  _T_132; 
  wire  _T_147; 
  wire  _T_149; 
  wire  _T_151; 
  wire  _T_152; 
  wire  _T_168; 
  wire  in_d_valid; 
  wire  _T_156; 
  wire [9:0] _GEN_17; 
  wire [9:0] _T_158; 
  wire  _T_162_1; 
  wire [2:0] da_bits_source; 
  wire [46:0] _T_186; 
  wire [46:0] _T_187; 
  dual_TLMonitor_4 dual_TLMonitor ( 
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_io_in_a_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt)
  );
  dual_Queue_2 a ( 
    .clock(a_clock),
    .reset(a_reset),
    .io_enq_ready(a_io_enq_ready),
    .io_enq_valid(a_io_enq_valid),
    .io_enq_bits_opcode(a_io_enq_bits_opcode),
    .io_enq_bits_size(a_io_enq_bits_size),
    .io_enq_bits_source(a_io_enq_bits_source),
    .io_deq_ready(a_io_deq_ready),
    .io_deq_valid(a_io_deq_valid),
    .io_deq_bits_opcode(a_io_deq_bits_opcode),
    .io_deq_bits_size(a_io_deq_bits_size),
    .io_deq_bits_source(a_io_deq_bits_source)
  );
  assign _T_6 = a_io_deq_ready & a_io_deq_valid; 
  assign _T_8 = 27'hfff << a_io_deq_bits_size; 
  assign _T_9 = _T_8[11:0]; 
  assign _T_10 = ~ _T_9; 
  assign _T_11 = _T_10[11:2]; 
  assign _T_12 = a_io_deq_bits_opcode[2]; 
  assign _T_13 = _T_12 == 1'h0; 
  assign _T_14 = _T_13 ? _T_11 : 10'h0; 
  assign _T_17 = _T_15 - 10'h1; 
  assign _T_18 = _T_15 == 10'h0; 
  assign _T_19 = _T_15 == 10'h1; 
  assign _T_20 = _T_14 == 10'h0; 
  assign a_last = _T_19 | _T_20; 
  assign _T_118 = _T_117 == 10'h0; 
  assign _T_50 = a_io_deq_valid & a_last; 
  assign da_valid = _T_50 & idle; 
  assign _T_120 = {da_valid,1'h0}; 
  assign _T_121 = {_T_120, 1'h0}; 
  assign _T_122 = _T_121[1:0]; 
  assign _T_123 = _T_120 | _T_122; 
  assign _T_125 = {_T_123, 1'h0}; 
  assign _T_126 = _T_125[1:0]; 
  assign _T_127 = ~ _T_126; 
  assign _T_129 = _T_127[1]; 
  assign _T_163_1 = _T_118 ? _T_129 : _T_161_1; 
  assign da_ready = auto_in_d_ready & _T_163_1; 
  assign _T_25 = da_ready & da_valid; 
  assign da_bits_size = a_io_deq_bits_size; 
  assign _T_27 = 27'hfff << da_bits_size; 
  assign _T_28 = _T_27[11:0]; 
  assign _T_29 = ~ _T_28; 
  assign _T_30 = _T_29[11:2]; 
  assign _GEN_4 = 3'h2 == a_io_deq_bits_opcode ? 3'h1 : 3'h0; 
  assign _GEN_5 = 3'h3 == a_io_deq_bits_opcode ? 3'h1 : _GEN_4; 
  assign _GEN_6 = 3'h4 == a_io_deq_bits_opcode ? 3'h1 : _GEN_5; 
  assign _GEN_7 = 3'h5 == a_io_deq_bits_opcode ? 3'h2 : _GEN_6; 
  assign _GEN_8 = 3'h6 == a_io_deq_bits_opcode ? 3'h4 : _GEN_7; 
  assign da_bits_opcode = 3'h7 == a_io_deq_bits_opcode ? 3'h4 : _GEN_8; 
  assign _T_31 = da_bits_opcode[0]; 
  assign _T_32 = _T_31 ? _T_30 : 10'h0; 
  assign _T_35 = _T_33 - 10'h1; 
  assign da_first = _T_33 == 10'h0; 
  assign _T_36 = _T_33 == 10'h1; 
  assign _T_37 = _T_32 == 10'h0; 
  assign da_last = _T_36 | _T_37; 
  assign _T_42 = idle | da_first; 
  assign _T_44 = _T_42 | reset; 
  assign _T_45 = _T_44 == 1'h0; 
  assign _T_46 = da_ready & da_last; 
  assign _T_47 = _T_46 & idle; 
  assign _T_48 = a_last == 1'h0; 
  assign _T_94 = da_bits_opcode == 3'h4; 
  assign _T_95 = _T_25 & _T_94; 
  assign _T_119 = _T_118 & auto_in_d_ready; 
  assign _T_132 = _T_129 & da_valid; 
  assign _T_147 = da_valid == 1'h0; 
  assign _T_149 = _T_147 | _T_132; 
  assign _T_151 = _T_149 | reset; 
  assign _T_152 = _T_151 == 1'h0; 
  assign _T_168 = _T_161_1 ? da_valid : 1'h0; 
  assign in_d_valid = _T_118 ? da_valid : _T_168; 
  assign _T_156 = auto_in_d_ready & in_d_valid; 
  assign _GEN_17 = {{9'd0}, _T_156}; 
  assign _T_158 = _T_117 - _GEN_17; 
  assign _T_162_1 = _T_118 ? _T_132 : _T_161_1; 
  assign da_bits_source = a_io_deq_bits_source; 
  assign _T_186 = {da_bits_opcode,2'h0,da_bits_size,da_bits_source,2'h1,32'h0,_T_31}; 
  assign _T_187 = _T_162_1 ? _T_186 : 47'h0; 
  assign auto_in_a_ready = a_io_enq_ready; 
  assign auto_in_d_valid = _T_118 ? da_valid : _T_168; 
  assign auto_in_d_bits_opcode = _T_187[46:44]; 
  assign auto_in_d_bits_param = _T_187[43:42]; 
  assign auto_in_d_bits_size = _T_187[41:38]; 
  assign auto_in_d_bits_source = _T_187[37:35]; 
  assign auto_in_d_bits_sink = _T_187[34]; 
  assign auto_in_d_bits_denied = _T_187[33]; 
  assign auto_in_d_bits_data = _T_187[32:1]; 
  assign auto_in_d_bits_corrupt = _T_187[0]; 
  assign TLMonitor_clock = clock; 
  assign TLMonitor_reset = reset; 
  assign TLMonitor_io_in_a_ready = a_io_enq_ready; 
  assign TLMonitor_io_in_a_valid = auto_in_a_valid; 
  assign TLMonitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; 
  assign TLMonitor_io_in_a_bits_param = auto_in_a_bits_param; 
  assign TLMonitor_io_in_a_bits_size = auto_in_a_bits_size; 
  assign TLMonitor_io_in_a_bits_source = auto_in_a_bits_source; 
  assign TLMonitor_io_in_a_bits_address = auto_in_a_bits_address; 
  assign TLMonitor_io_in_a_bits_mask = auto_in_a_bits_mask; 
  assign TLMonitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; 
  assign TLMonitor_io_in_d_ready = auto_in_d_ready; 
  assign TLMonitor_io_in_d_valid = _T_118 ? da_valid : _T_168; 
  assign TLMonitor_io_in_d_bits_opcode = _T_187[46:44]; 
  assign TLMonitor_io_in_d_bits_param = _T_187[43:42]; 
  assign TLMonitor_io_in_d_bits_size = _T_187[41:38]; 
  assign TLMonitor_io_in_d_bits_source = _T_187[37:35]; 
  assign TLMonitor_io_in_d_bits_sink = _T_187[34]; 
  assign TLMonitor_io_in_d_bits_denied = _T_187[33]; 
  assign TLMonitor_io_in_d_bits_corrupt = _T_187[0]; 
  assign a_clock = clock; 
  assign a_reset = reset; 
  assign a_io_enq_valid = auto_in_a_valid; 
  assign a_io_enq_bits_opcode = auto_in_a_bits_opcode; 
  assign a_io_enq_bits_size = auto_in_a_bits_size; 
  assign a_io_enq_bits_source = auto_in_a_bits_source; 
  assign a_io_deq_ready = _T_47 | _T_48; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  idle = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_15 = _RAND_1[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_117 = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_161_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_33 = _RAND_4[9:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      idle <= 1'h1;
    end else begin
      if (_T_95) begin
        idle <= 1'h0;
      end
    end
    if (reset) begin
      _T_15 <= 10'h0;
    end else begin
      if (_T_6) begin
        if (_T_18) begin
          if (_T_13) begin
            _T_15 <= _T_11;
          end else begin
            _T_15 <= 10'h0;
          end
        end else begin
          _T_15 <= _T_17;
        end
      end
    end
    if (reset) begin
      _T_117 <= 10'h0;
    end else begin
      if (_T_119) begin
        if (_T_132) begin
          if (_T_31) begin
            _T_117 <= _T_30;
          end else begin
            _T_117 <= 10'h0;
          end
        end else begin
          _T_117 <= 10'h0;
        end
      end else begin
        _T_117 <= _T_158;
      end
    end
    if (reset) begin
      _T_161_1 <= 1'h0;
    end else begin
      if (_T_118) begin
        _T_161_1 <= _T_132;
      end
    end
    if (reset) begin
      _T_33 <= 10'h0;
    end else begin
      if (_T_25) begin
        if (da_first) begin
          if (_T_31) begin
            _T_33 <= _T_30;
          end else begin
            _T_33 <= 10'h0;
          end
        end else begin
          _T_33 <= _T_35;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_45) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Error.scala:28 assert (idle || da_first) // we only send Grant, never GrantData => simplified flow control below\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_45) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_152) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:70 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_152) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLError_2( 
  input         clock, 
  input         reset, 
  output        auto_in_a_ready, 
  input         auto_in_a_valid, 
  input  [2:0]  auto_in_a_bits_opcode, 
  input  [2:0]  auto_in_a_bits_param, 
  input  [2:0]  auto_in_a_bits_size, 
  input  [6:0]  auto_in_a_bits_source, 
  input  [28:0] auto_in_a_bits_address, 
  input  [3:0]  auto_in_a_bits_mask, 
  input         auto_in_a_bits_corrupt, 
  output        auto_in_c_ready, 
  input         auto_in_c_valid, 
  input  [2:0]  auto_in_c_bits_opcode, 
  input  [2:0]  auto_in_c_bits_param, 
  input  [2:0]  auto_in_c_bits_size, 
  input  [6:0]  auto_in_c_bits_source, 
  input  [28:0] auto_in_c_bits_address, 
  input         auto_in_c_bits_corrupt, 
  input         auto_in_d_ready, 
  output        auto_in_d_valid, 
  output [2:0]  auto_in_d_bits_opcode, 
  output [1:0]  auto_in_d_bits_param, 
  output [2:0]  auto_in_d_bits_size, 
  output [6:0]  auto_in_d_bits_source, 
  output        auto_in_d_bits_sink, 
  output        auto_in_d_bits_denied, 
  output [31:0] auto_in_d_bits_data, 
  output        auto_in_d_bits_corrupt, 
  input         auto_in_e_valid 
);
  wire  TLMonitor_clock; 
  wire  TLMonitor_reset; 
  wire  TLMonitor_io_in_a_ready; 
  wire  TLMonitor_io_in_a_valid; 
  wire [2:0] TLMonitor_io_in_a_bits_opcode; 
  wire [2:0] TLMonitor_io_in_a_bits_param; 
  wire [2:0] TLMonitor_io_in_a_bits_size; 
  wire [6:0] TLMonitor_io_in_a_bits_source; 
  wire [28:0] TLMonitor_io_in_a_bits_address; 
  wire [3:0] TLMonitor_io_in_a_bits_mask; 
  wire  TLMonitor_io_in_a_bits_corrupt; 
  wire  TLMonitor_io_in_c_ready; 
  wire  TLMonitor_io_in_c_valid; 
  wire [2:0] TLMonitor_io_in_c_bits_opcode; 
  wire [2:0] TLMonitor_io_in_c_bits_param; 
  wire [2:0] TLMonitor_io_in_c_bits_size; 
  wire [6:0] TLMonitor_io_in_c_bits_source; 
  wire [28:0] TLMonitor_io_in_c_bits_address; 
  wire  TLMonitor_io_in_c_bits_corrupt; 
  wire  TLMonitor_io_in_d_ready; 
  wire  TLMonitor_io_in_d_valid; 
  wire [2:0] TLMonitor_io_in_d_bits_opcode; 
  wire [1:0] TLMonitor_io_in_d_bits_param; 
  wire [2:0] TLMonitor_io_in_d_bits_size; 
  wire [6:0] TLMonitor_io_in_d_bits_source; 
  wire  TLMonitor_io_in_d_bits_sink; 
  wire  TLMonitor_io_in_d_bits_denied; 
  wire  TLMonitor_io_in_d_bits_corrupt; 
  wire  TLMonitor_io_in_e_valid; 
  wire  a_clock; 
  wire  a_reset; 
  wire  a_io_enq_ready; 
  wire  a_io_enq_valid; 
  wire [2:0] a_io_enq_bits_opcode; 
  wire [2:0] a_io_enq_bits_size; 
  wire [6:0] a_io_enq_bits_source; 
  wire  a_io_deq_ready; 
  wire  a_io_deq_valid; 
  wire [2:0] a_io_deq_bits_opcode; 
  wire [2:0] a_io_deq_bits_size; 
  wire [6:0] a_io_deq_bits_source; 
  wire  Queue_clock; 
  wire  Queue_reset; 
  wire  Queue_io_enq_ready; 
  wire  Queue_io_enq_valid; 
  wire [2:0] Queue_io_enq_bits_opcode; 
  wire [2:0] Queue_io_enq_bits_param; 
  wire [2:0] Queue_io_enq_bits_size; 
  wire [6:0] Queue_io_enq_bits_source; 
  wire  Queue_io_deq_ready; 
  wire  Queue_io_deq_valid; 
  wire [2:0] Queue_io_deq_bits_opcode; 
  wire [2:0] Queue_io_deq_bits_param; 
  wire [2:0] Queue_io_deq_bits_size; 
  wire [6:0] Queue_io_deq_bits_source; 
  reg  idle; 
  reg [31:0] _RAND_0;
  wire  _T_6; 
  wire [12:0] _T_8; 
  wire [5:0] _T_9; 
  wire [5:0] _T_10; 
  wire [3:0] _T_11; 
  wire  _T_12; 
  wire  _T_13; 
  wire [3:0] _T_14; 
  reg [3:0] _T_15; 
  reg [31:0] _RAND_1;
  wire [3:0] _T_17; 
  wire  _T_18; 
  wire  _T_19; 
  wire  _T_20; 
  wire  a_last; 
  reg [3:0] _T_117; 
  reg [31:0] _RAND_2;
  wire  _T_118; 
  wire  _T_50; 
  wire  da_valid; 
  reg [3:0] _T_63; 
  reg [31:0] _RAND_3;
  wire  _T_67; 
  wire  _T_61; 
  wire [12:0] _T_57; 
  wire [5:0] _T_58; 
  wire [5:0] _T_59; 
  wire [3:0] _T_60; 
  wire [3:0] _T_62; 
  wire  _T_68; 
  wire  _T_69; 
  wire  _T_100; 
  wire [1:0] _T_120; 
  wire [2:0] _T_121; 
  wire [1:0] _T_122; 
  wire [1:0] _T_123; 
  wire [2:0] _T_125; 
  wire [1:0] _T_126; 
  wire [1:0] _T_127; 
  wire  _T_129; 
  reg  _T_161_1; 
  reg [31:0] _RAND_4;
  wire  _T_163_1; 
  wire  da_ready; 
  wire  _T_25; 
  wire [2:0] da_bits_size; 
  wire [12:0] _T_27; 
  wire [5:0] _T_28; 
  wire [5:0] _T_29; 
  wire [3:0] _T_30; 
  wire [2:0] _GEN_4; 
  wire [2:0] _GEN_5; 
  wire [2:0] _GEN_6; 
  wire [2:0] _GEN_7; 
  wire [2:0] _GEN_8; 
  wire [2:0] da_bits_opcode; 
  wire  _T_31; 
  wire [3:0] _T_32; 
  reg [3:0] _T_33; 
  reg [31:0] _RAND_5;
  wire [3:0] _T_35; 
  wire  da_first; 
  wire  _T_36; 
  wire  _T_37; 
  wire  da_last; 
  wire  _T_42; 
  wire  _T_44; 
  wire  _T_45; 
  wire  _T_46; 
  wire  _T_47; 
  wire  _T_48; 
  wire  _T_55; 
  wire [3:0] _T_65; 
  wire  _T_66; 
  wire  _T_128; 
  reg  _T_161_0; 
  reg [31:0] _RAND_6;
  wire  _T_163_0; 
  wire  _T_164; 
  wire [2:0] _T_54_bits_size; 
  wire  _T_94; 
  wire  _T_95; 
  wire  _T_98; 
  wire [1:0] _T_102; 
  wire [1:0] _GEN_15; 
  wire [1:0] _GEN_16; 
  wire  _T_119; 
  wire  _T_131; 
  wire  _T_132; 
  wire  _T_135; 
  wire  _T_137; 
  wire  _T_140; 
  wire  _T_141; 
  wire  _T_144; 
  wire  _T_145; 
  wire  _T_146; 
  wire  _T_147; 
  wire  _T_149; 
  wire  _T_151; 
  wire  _T_152; 
  wire  _T_167; 
  wire  _T_168; 
  wire  _T_169; 
  wire  in_d_valid; 
  wire  _T_156; 
  wire [3:0] _GEN_17; 
  wire [3:0] _T_158; 
  wire  _T_162_0; 
  wire  _T_162_1; 
  wire [6:0] _T_54_bits_source; 
  wire [49:0] _T_178; 
  wire [49:0] _T_179; 
  wire [6:0] da_bits_source; 
  wire [49:0] _T_186; 
  wire [49:0] _T_187; 
  wire [49:0] _T_188; 
  dual_TLMonitor_13 dual_TLMonitor ( 
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_io_in_a_bits_corrupt),
    .io_in_c_ready(TLMonitor_io_in_c_ready),
    .io_in_c_valid(TLMonitor_io_in_c_valid),
    .io_in_c_bits_opcode(TLMonitor_io_in_c_bits_opcode),
    .io_in_c_bits_param(TLMonitor_io_in_c_bits_param),
    .io_in_c_bits_size(TLMonitor_io_in_c_bits_size),
    .io_in_c_bits_source(TLMonitor_io_in_c_bits_source),
    .io_in_c_bits_address(TLMonitor_io_in_c_bits_address),
    .io_in_c_bits_corrupt(TLMonitor_io_in_c_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt),
    .io_in_e_valid(TLMonitor_io_in_e_valid)
  );
  dual_Queue_67 a ( 
    .clock(a_clock),
    .reset(a_reset),
    .io_enq_ready(a_io_enq_ready),
    .io_enq_valid(a_io_enq_valid),
    .io_enq_bits_opcode(a_io_enq_bits_opcode),
    .io_enq_bits_size(a_io_enq_bits_size),
    .io_enq_bits_source(a_io_enq_bits_source),
    .io_deq_ready(a_io_deq_ready),
    .io_deq_valid(a_io_deq_valid),
    .io_deq_bits_opcode(a_io_deq_bits_opcode),
    .io_deq_bits_size(a_io_deq_bits_size),
    .io_deq_bits_source(a_io_deq_bits_source)
  );
  dual_Queue_68 dual_Queue ( 
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_opcode(Queue_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_io_enq_bits_param),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_source(Queue_io_enq_bits_source),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_opcode(Queue_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_io_deq_bits_param),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_source(Queue_io_deq_bits_source)
  );
  assign _T_6 = a_io_deq_ready & a_io_deq_valid; 
  assign _T_8 = 13'h3f << a_io_deq_bits_size; 
  assign _T_9 = _T_8[5:0]; 
  assign _T_10 = ~ _T_9; 
  assign _T_11 = _T_10[5:2]; 
  assign _T_12 = a_io_deq_bits_opcode[2]; 
  assign _T_13 = _T_12 == 1'h0; 
  assign _T_14 = _T_13 ? _T_11 : 4'h0; 
  assign _T_17 = _T_15 - 4'h1; 
  assign _T_18 = _T_15 == 4'h0; 
  assign _T_19 = _T_15 == 4'h1; 
  assign _T_20 = _T_14 == 4'h0; 
  assign a_last = _T_19 | _T_20; 
  assign _T_118 = _T_117 == 4'h0; 
  assign _T_50 = a_io_deq_valid & a_last; 
  assign da_valid = _T_50 & idle; 
  assign _T_67 = _T_63 == 4'h1; 
  assign _T_61 = Queue_io_deq_bits_opcode[0]; 
  assign _T_57 = 13'h3f << Queue_io_deq_bits_size; 
  assign _T_58 = _T_57[5:0]; 
  assign _T_59 = ~ _T_58; 
  assign _T_60 = _T_59[5:2]; 
  assign _T_62 = _T_61 ? _T_60 : 4'h0; 
  assign _T_68 = _T_62 == 4'h0; 
  assign _T_69 = _T_67 | _T_68; 
  assign _T_100 = Queue_io_deq_valid & _T_69; 
  assign _T_120 = {da_valid,_T_100}; 
  assign _T_121 = {_T_120, 1'h0}; 
  assign _T_122 = _T_121[1:0]; 
  assign _T_123 = _T_120 | _T_122; 
  assign _T_125 = {_T_123, 1'h0}; 
  assign _T_126 = _T_125[1:0]; 
  assign _T_127 = ~ _T_126; 
  assign _T_129 = _T_127[1]; 
  assign _T_163_1 = _T_118 ? _T_129 : _T_161_1; 
  assign da_ready = auto_in_d_ready & _T_163_1; 
  assign _T_25 = da_ready & da_valid; 
  assign da_bits_size = a_io_deq_bits_size; 
  assign _T_27 = 13'h3f << da_bits_size; 
  assign _T_28 = _T_27[5:0]; 
  assign _T_29 = ~ _T_28; 
  assign _T_30 = _T_29[5:2]; 
  assign _GEN_4 = 3'h2 == a_io_deq_bits_opcode ? 3'h1 : 3'h0; 
  assign _GEN_5 = 3'h3 == a_io_deq_bits_opcode ? 3'h1 : _GEN_4; 
  assign _GEN_6 = 3'h4 == a_io_deq_bits_opcode ? 3'h1 : _GEN_5; 
  assign _GEN_7 = 3'h5 == a_io_deq_bits_opcode ? 3'h2 : _GEN_6; 
  assign _GEN_8 = 3'h6 == a_io_deq_bits_opcode ? 3'h4 : _GEN_7; 
  assign da_bits_opcode = 3'h7 == a_io_deq_bits_opcode ? 3'h4 : _GEN_8; 
  assign _T_31 = da_bits_opcode[0]; 
  assign _T_32 = _T_31 ? _T_30 : 4'h0; 
  assign _T_35 = _T_33 - 4'h1; 
  assign da_first = _T_33 == 4'h0; 
  assign _T_36 = _T_33 == 4'h1; 
  assign _T_37 = _T_32 == 4'h0; 
  assign da_last = _T_36 | _T_37; 
  assign _T_42 = idle | da_first; 
  assign _T_44 = _T_42 | reset; 
  assign _T_45 = _T_44 == 1'h0; 
  assign _T_46 = da_ready & da_last; 
  assign _T_47 = _T_46 & idle; 
  assign _T_48 = a_last == 1'h0; 
  assign _T_55 = Queue_io_deq_ready & Queue_io_deq_valid; 
  assign _T_65 = _T_63 - 4'h1; 
  assign _T_66 = _T_63 == 4'h0; 
  assign _T_128 = _T_127[0]; 
  assign _T_163_0 = _T_118 ? _T_128 : _T_161_0; 
  assign _T_164 = auto_in_d_ready & _T_163_0; 
  assign _T_54_bits_size = Queue_io_deq_bits_size; 
  assign _T_94 = da_bits_opcode == 3'h4; 
  assign _T_95 = _T_25 & _T_94; 
  assign _T_98 = _T_69 == 1'h0; 
  assign _T_102 = Queue_io_deq_bits_param[1:0]; 
  assign _GEN_15 = 2'h1 == _T_102 ? 2'h2 : 2'h1; 
  assign _GEN_16 = 2'h2 == _T_102 ? 2'h2 : _GEN_15; 
  assign _T_119 = _T_118 & auto_in_d_ready; 
  assign _T_131 = _T_128 & _T_100; 
  assign _T_132 = _T_129 & da_valid; 
  assign _T_135 = _T_131 | _T_132; 
  assign _T_137 = _T_131 == 1'h0; 
  assign _T_140 = _T_132 == 1'h0; 
  assign _T_141 = _T_137 | _T_140; 
  assign _T_144 = _T_141 | reset; 
  assign _T_145 = _T_144 == 1'h0; 
  assign _T_146 = _T_100 | da_valid; 
  assign _T_147 = _T_146 == 1'h0; 
  assign _T_149 = _T_147 | _T_135; 
  assign _T_151 = _T_149 | reset; 
  assign _T_152 = _T_151 == 1'h0; 
  assign _T_167 = _T_161_0 ? _T_100 : 1'h0; 
  assign _T_168 = _T_161_1 ? da_valid : 1'h0; 
  assign _T_169 = _T_167 | _T_168; 
  assign in_d_valid = _T_118 ? _T_146 : _T_169; 
  assign _T_156 = auto_in_d_ready & in_d_valid; 
  assign _GEN_17 = {{3'd0}, _T_156}; 
  assign _T_158 = _T_117 - _GEN_17; 
  assign _T_162_0 = _T_118 ? _T_131 : _T_161_0; 
  assign _T_162_1 = _T_118 ? _T_132 : _T_161_1; 
  assign _T_54_bits_source = Queue_io_deq_bits_source; 
  assign _T_178 = {3'h6,_GEN_16,_T_54_bits_size,_T_54_bits_source,35'h0}; 
  assign _T_179 = _T_162_0 ? _T_178 : 50'h0; 
  assign da_bits_source = a_io_deq_bits_source; 
  assign _T_186 = {da_bits_opcode,2'h0,da_bits_size,da_bits_source,2'h1,32'h0,_T_31}; 
  assign _T_187 = _T_162_1 ? _T_186 : 50'h0; 
  assign _T_188 = _T_179 | _T_187; 
  assign auto_in_a_ready = a_io_enq_ready; 
  assign auto_in_c_ready = Queue_io_enq_ready; 
  assign auto_in_d_valid = _T_118 ? _T_146 : _T_169; 
  assign auto_in_d_bits_opcode = _T_188[49:47]; 
  assign auto_in_d_bits_param = _T_188[46:45]; 
  assign auto_in_d_bits_size = _T_188[44:42]; 
  assign auto_in_d_bits_source = _T_188[41:35]; 
  assign auto_in_d_bits_sink = _T_188[34]; 
  assign auto_in_d_bits_denied = _T_188[33]; 
  assign auto_in_d_bits_data = _T_188[32:1]; 
  assign auto_in_d_bits_corrupt = _T_188[0]; 
  assign TLMonitor_clock = clock; 
  assign TLMonitor_reset = reset; 
  assign TLMonitor_io_in_a_ready = a_io_enq_ready; 
  assign TLMonitor_io_in_a_valid = auto_in_a_valid; 
  assign TLMonitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; 
  assign TLMonitor_io_in_a_bits_param = auto_in_a_bits_param; 
  assign TLMonitor_io_in_a_bits_size = auto_in_a_bits_size; 
  assign TLMonitor_io_in_a_bits_source = auto_in_a_bits_source; 
  assign TLMonitor_io_in_a_bits_address = auto_in_a_bits_address; 
  assign TLMonitor_io_in_a_bits_mask = auto_in_a_bits_mask; 
  assign TLMonitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; 
  assign TLMonitor_io_in_c_ready = Queue_io_enq_ready; 
  assign TLMonitor_io_in_c_valid = auto_in_c_valid; 
  assign TLMonitor_io_in_c_bits_opcode = auto_in_c_bits_opcode; 
  assign TLMonitor_io_in_c_bits_param = auto_in_c_bits_param; 
  assign TLMonitor_io_in_c_bits_size = auto_in_c_bits_size; 
  assign TLMonitor_io_in_c_bits_source = auto_in_c_bits_source; 
  assign TLMonitor_io_in_c_bits_address = auto_in_c_bits_address; 
  assign TLMonitor_io_in_c_bits_corrupt = auto_in_c_bits_corrupt; 
  assign TLMonitor_io_in_d_ready = auto_in_d_ready; 
  assign TLMonitor_io_in_d_valid = _T_118 ? _T_146 : _T_169; 
  assign TLMonitor_io_in_d_bits_opcode = _T_188[49:47]; 
  assign TLMonitor_io_in_d_bits_param = _T_188[46:45]; 
  assign TLMonitor_io_in_d_bits_size = _T_188[44:42]; 
  assign TLMonitor_io_in_d_bits_source = _T_188[41:35]; 
  assign TLMonitor_io_in_d_bits_sink = _T_188[34]; 
  assign TLMonitor_io_in_d_bits_denied = _T_188[33]; 
  assign TLMonitor_io_in_d_bits_corrupt = _T_188[0]; 
  assign TLMonitor_io_in_e_valid = auto_in_e_valid; 
  assign a_clock = clock; 
  assign a_reset = reset; 
  assign a_io_enq_valid = auto_in_a_valid; 
  assign a_io_enq_bits_opcode = auto_in_a_bits_opcode; 
  assign a_io_enq_bits_size = auto_in_a_bits_size; 
  assign a_io_enq_bits_source = auto_in_a_bits_source; 
  assign a_io_deq_ready = _T_47 | _T_48; 
  assign Queue_clock = clock; 
  assign Queue_reset = reset; 
  assign Queue_io_enq_valid = auto_in_c_valid; 
  assign Queue_io_enq_bits_opcode = auto_in_c_bits_opcode; 
  assign Queue_io_enq_bits_param = auto_in_c_bits_param; 
  assign Queue_io_enq_bits_size = auto_in_c_bits_size; 
  assign Queue_io_enq_bits_source = auto_in_c_bits_source; 
  assign Queue_io_deq_ready = _T_164 | _T_98; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  idle = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_15 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_117 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_63 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_161_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_33 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_161_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      idle <= 1'h1;
    end else begin
      if (auto_in_e_valid) begin
        idle <= 1'h1;
      end else begin
        if (_T_95) begin
          idle <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_15 <= 4'h0;
    end else begin
      if (_T_6) begin
        if (_T_18) begin
          if (_T_13) begin
            _T_15 <= _T_11;
          end else begin
            _T_15 <= 4'h0;
          end
        end else begin
          _T_15 <= _T_17;
        end
      end
    end
    if (reset) begin
      _T_117 <= 4'h0;
    end else begin
      if (_T_119) begin
        if (_T_132) begin
          if (_T_31) begin
            _T_117 <= _T_30;
          end else begin
            _T_117 <= 4'h0;
          end
        end else begin
          _T_117 <= 4'h0;
        end
      end else begin
        _T_117 <= _T_158;
      end
    end
    if (reset) begin
      _T_63 <= 4'h0;
    end else begin
      if (_T_55) begin
        if (_T_66) begin
          if (_T_61) begin
            _T_63 <= _T_60;
          end else begin
            _T_63 <= 4'h0;
          end
        end else begin
          _T_63 <= _T_65;
        end
      end
    end
    if (reset) begin
      _T_161_1 <= 1'h0;
    end else begin
      if (_T_118) begin
        _T_161_1 <= _T_132;
      end
    end
    if (reset) begin
      _T_33 <= 4'h0;
    end else begin
      if (_T_25) begin
        if (da_first) begin
          if (_T_31) begin
            _T_33 <= _T_30;
          end else begin
            _T_33 <= 4'h0;
          end
        end else begin
          _T_33 <= _T_35;
        end
      end
    end
    if (reset) begin
      _T_161_0 <= 1'h0;
    end else begin
      if (_T_118) begin
        _T_161_0 <= _T_131;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_45) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Error.scala:28 assert (idle || da_first) // we only send Grant, never GrantData => simplified flow control below\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_45) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_145) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_145) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_152) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:70 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_152) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLError( 
  input         clock, 
  input         reset, 
  output        auto_in_a_ready, 
  input         auto_in_a_valid, 
  input  [2:0]  auto_in_a_bits_opcode, 
  input  [2:0]  auto_in_a_bits_param, 
  input  [2:0]  auto_in_a_bits_size, 
  input  [2:0]  auto_in_a_bits_source, 
  input  [28:0] auto_in_a_bits_address, 
  input  [3:0]  auto_in_a_bits_mask, 
  input         auto_in_a_bits_corrupt, 
  input         auto_in_d_ready, 
  output        auto_in_d_valid, 
  output [2:0]  auto_in_d_bits_opcode, 
  output [1:0]  auto_in_d_bits_param, 
  output [2:0]  auto_in_d_bits_size, 
  output [2:0]  auto_in_d_bits_source, 
  output        auto_in_d_bits_sink, 
  output        auto_in_d_bits_denied, 
  output [31:0] auto_in_d_bits_data, 
  output        auto_in_d_bits_corrupt 
);
  wire  TLMonitor_clock; 
  wire  TLMonitor_reset; 
  wire  TLMonitor_io_in_a_ready; 
  wire  TLMonitor_io_in_a_valid; 
  wire [2:0] TLMonitor_io_in_a_bits_opcode; 
  wire [2:0] TLMonitor_io_in_a_bits_param; 
  wire [2:0] TLMonitor_io_in_a_bits_size; 
  wire [2:0] TLMonitor_io_in_a_bits_source; 
  wire [28:0] TLMonitor_io_in_a_bits_address; 
  wire [3:0] TLMonitor_io_in_a_bits_mask; 
  wire  TLMonitor_io_in_a_bits_corrupt; 
  wire  TLMonitor_io_in_d_ready; 
  wire  TLMonitor_io_in_d_valid; 
  wire [2:0] TLMonitor_io_in_d_bits_opcode; 
  wire [1:0] TLMonitor_io_in_d_bits_param; 
  wire [2:0] TLMonitor_io_in_d_bits_size; 
  wire [2:0] TLMonitor_io_in_d_bits_source; 
  wire  TLMonitor_io_in_d_bits_sink; 
  wire  TLMonitor_io_in_d_bits_denied; 
  wire  TLMonitor_io_in_d_bits_corrupt; 
  wire  a_clock; 
  wire  a_reset; 
  wire  a_io_enq_ready; 
  wire  a_io_enq_valid; 
  wire [2:0] a_io_enq_bits_opcode; 
  wire [2:0] a_io_enq_bits_size; 
  wire [2:0] a_io_enq_bits_source; 
  wire  a_io_deq_ready; 
  wire  a_io_deq_valid; 
  wire [2:0] a_io_deq_bits_opcode; 
  wire [2:0] a_io_deq_bits_size; 
  wire [2:0] a_io_deq_bits_source; 
  reg  idle; 
  reg [31:0] _RAND_0;
  wire  _T_6; 
  wire [12:0] _T_8; 
  wire [5:0] _T_9; 
  wire [5:0] _T_10; 
  wire [3:0] _T_11; 
  wire  _T_12; 
  wire  _T_13; 
  wire [3:0] _T_14; 
  reg [3:0] _T_15; 
  reg [31:0] _RAND_1;
  wire [3:0] _T_17; 
  wire  _T_18; 
  wire  _T_19; 
  wire  _T_20; 
  wire  a_last; 
  reg [3:0] _T_117; 
  reg [31:0] _RAND_2;
  wire  _T_118; 
  wire  _T_50; 
  wire  da_valid; 
  wire [1:0] _T_120; 
  wire [2:0] _T_121; 
  wire [1:0] _T_122; 
  wire [1:0] _T_123; 
  wire [2:0] _T_125; 
  wire [1:0] _T_126; 
  wire [1:0] _T_127; 
  wire  _T_129; 
  reg  _T_161_1; 
  reg [31:0] _RAND_3;
  wire  _T_163_1; 
  wire  da_ready; 
  wire  _T_25; 
  wire [2:0] da_bits_size; 
  wire [12:0] _T_27; 
  wire [5:0] _T_28; 
  wire [5:0] _T_29; 
  wire [3:0] _T_30; 
  wire [2:0] _GEN_4; 
  wire [2:0] _GEN_5; 
  wire [2:0] _GEN_6; 
  wire [2:0] _GEN_7; 
  wire [2:0] _GEN_8; 
  wire [2:0] da_bits_opcode; 
  wire  _T_31; 
  wire [3:0] _T_32; 
  reg [3:0] _T_33; 
  reg [31:0] _RAND_4;
  wire [3:0] _T_35; 
  wire  da_first; 
  wire  _T_36; 
  wire  _T_37; 
  wire  da_last; 
  wire  _T_42; 
  wire  _T_44; 
  wire  _T_45; 
  wire  _T_46; 
  wire  _T_47; 
  wire  _T_48; 
  wire  _T_94; 
  wire  _T_95; 
  wire  _T_119; 
  wire  _T_132; 
  wire  _T_147; 
  wire  _T_149; 
  wire  _T_151; 
  wire  _T_152; 
  wire  _T_168; 
  wire  in_d_valid; 
  wire  _T_156; 
  wire [3:0] _GEN_17; 
  wire [3:0] _T_158; 
  wire  _T_162_1; 
  wire [2:0] da_bits_source; 
  wire [45:0] _T_186; 
  wire [45:0] _T_187; 
  dual_TLMonitor_2 dual_TLMonitor ( 
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_io_in_a_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt)
  );
  dual_Queue a ( 
    .clock(a_clock),
    .reset(a_reset),
    .io_enq_ready(a_io_enq_ready),
    .io_enq_valid(a_io_enq_valid),
    .io_enq_bits_opcode(a_io_enq_bits_opcode),
    .io_enq_bits_size(a_io_enq_bits_size),
    .io_enq_bits_source(a_io_enq_bits_source),
    .io_deq_ready(a_io_deq_ready),
    .io_deq_valid(a_io_deq_valid),
    .io_deq_bits_opcode(a_io_deq_bits_opcode),
    .io_deq_bits_size(a_io_deq_bits_size),
    .io_deq_bits_source(a_io_deq_bits_source)
  );
  assign _T_6 = a_io_deq_ready & a_io_deq_valid; 
  assign _T_8 = 13'h3f << a_io_deq_bits_size; 
  assign _T_9 = _T_8[5:0]; 
  assign _T_10 = ~ _T_9; 
  assign _T_11 = _T_10[5:2]; 
  assign _T_12 = a_io_deq_bits_opcode[2]; 
  assign _T_13 = _T_12 == 1'h0; 
  assign _T_14 = _T_13 ? _T_11 : 4'h0; 
  assign _T_17 = _T_15 - 4'h1; 
  assign _T_18 = _T_15 == 4'h0; 
  assign _T_19 = _T_15 == 4'h1; 
  assign _T_20 = _T_14 == 4'h0; 
  assign a_last = _T_19 | _T_20; 
  assign _T_118 = _T_117 == 4'h0; 
  assign _T_50 = a_io_deq_valid & a_last; 
  assign da_valid = _T_50 & idle; 
  assign _T_120 = {da_valid,1'h0}; 
  assign _T_121 = {_T_120, 1'h0}; 
  assign _T_122 = _T_121[1:0]; 
  assign _T_123 = _T_120 | _T_122; 
  assign _T_125 = {_T_123, 1'h0}; 
  assign _T_126 = _T_125[1:0]; 
  assign _T_127 = ~ _T_126; 
  assign _T_129 = _T_127[1]; 
  assign _T_163_1 = _T_118 ? _T_129 : _T_161_1; 
  assign da_ready = auto_in_d_ready & _T_163_1; 
  assign _T_25 = da_ready & da_valid; 
  assign da_bits_size = a_io_deq_bits_size; 
  assign _T_27 = 13'h3f << da_bits_size; 
  assign _T_28 = _T_27[5:0]; 
  assign _T_29 = ~ _T_28; 
  assign _T_30 = _T_29[5:2]; 
  assign _GEN_4 = 3'h2 == a_io_deq_bits_opcode ? 3'h1 : 3'h0; 
  assign _GEN_5 = 3'h3 == a_io_deq_bits_opcode ? 3'h1 : _GEN_4; 
  assign _GEN_6 = 3'h4 == a_io_deq_bits_opcode ? 3'h1 : _GEN_5; 
  assign _GEN_7 = 3'h5 == a_io_deq_bits_opcode ? 3'h2 : _GEN_6; 
  assign _GEN_8 = 3'h6 == a_io_deq_bits_opcode ? 3'h4 : _GEN_7; 
  assign da_bits_opcode = 3'h7 == a_io_deq_bits_opcode ? 3'h4 : _GEN_8; 
  assign _T_31 = da_bits_opcode[0]; 
  assign _T_32 = _T_31 ? _T_30 : 4'h0; 
  assign _T_35 = _T_33 - 4'h1; 
  assign da_first = _T_33 == 4'h0; 
  assign _T_36 = _T_33 == 4'h1; 
  assign _T_37 = _T_32 == 4'h0; 
  assign da_last = _T_36 | _T_37; 
  assign _T_42 = idle | da_first; 
  assign _T_44 = _T_42 | reset; 
  assign _T_45 = _T_44 == 1'h0; 
  assign _T_46 = da_ready & da_last; 
  assign _T_47 = _T_46 & idle; 
  assign _T_48 = a_last == 1'h0; 
  assign _T_94 = da_bits_opcode == 3'h4; 
  assign _T_95 = _T_25 & _T_94; 
  assign _T_119 = _T_118 & auto_in_d_ready; 
  assign _T_132 = _T_129 & da_valid; 
  assign _T_147 = da_valid == 1'h0; 
  assign _T_149 = _T_147 | _T_132; 
  assign _T_151 = _T_149 | reset; 
  assign _T_152 = _T_151 == 1'h0; 
  assign _T_168 = _T_161_1 ? da_valid : 1'h0; 
  assign in_d_valid = _T_118 ? da_valid : _T_168; 
  assign _T_156 = auto_in_d_ready & in_d_valid; 
  assign _GEN_17 = {{3'd0}, _T_156}; 
  assign _T_158 = _T_117 - _GEN_17; 
  assign _T_162_1 = _T_118 ? _T_132 : _T_161_1; 
  assign da_bits_source = a_io_deq_bits_source; 
  assign _T_186 = {da_bits_opcode,2'h0,da_bits_size,da_bits_source,2'h1,32'h0,_T_31}; 
  assign _T_187 = _T_162_1 ? _T_186 : 46'h0; 
  assign auto_in_a_ready = a_io_enq_ready; 
  assign auto_in_d_valid = _T_118 ? da_valid : _T_168; 
  assign auto_in_d_bits_opcode = _T_187[45:43]; 
  assign auto_in_d_bits_param = _T_187[42:41]; 
  assign auto_in_d_bits_size = _T_187[40:38]; 
  assign auto_in_d_bits_source = _T_187[37:35]; 
  assign auto_in_d_bits_sink = _T_187[34]; 
  assign auto_in_d_bits_denied = _T_187[33]; 
  assign auto_in_d_bits_data = _T_187[32:1]; 
  assign auto_in_d_bits_corrupt = _T_187[0]; 
  assign TLMonitor_clock = clock; 
  assign TLMonitor_reset = reset; 
  assign TLMonitor_io_in_a_ready = a_io_enq_ready; 
  assign TLMonitor_io_in_a_valid = auto_in_a_valid; 
  assign TLMonitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; 
  assign TLMonitor_io_in_a_bits_param = auto_in_a_bits_param; 
  assign TLMonitor_io_in_a_bits_size = auto_in_a_bits_size; 
  assign TLMonitor_io_in_a_bits_source = auto_in_a_bits_source; 
  assign TLMonitor_io_in_a_bits_address = auto_in_a_bits_address; 
  assign TLMonitor_io_in_a_bits_mask = auto_in_a_bits_mask; 
  assign TLMonitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; 
  assign TLMonitor_io_in_d_ready = auto_in_d_ready; 
  assign TLMonitor_io_in_d_valid = _T_118 ? da_valid : _T_168; 
  assign TLMonitor_io_in_d_bits_opcode = _T_187[45:43]; 
  assign TLMonitor_io_in_d_bits_param = _T_187[42:41]; 
  assign TLMonitor_io_in_d_bits_size = _T_187[40:38]; 
  assign TLMonitor_io_in_d_bits_source = _T_187[37:35]; 
  assign TLMonitor_io_in_d_bits_sink = _T_187[34]; 
  assign TLMonitor_io_in_d_bits_denied = _T_187[33]; 
  assign TLMonitor_io_in_d_bits_corrupt = _T_187[0]; 
  assign a_clock = clock; 
  assign a_reset = reset; 
  assign a_io_enq_valid = auto_in_a_valid; 
  assign a_io_enq_bits_opcode = auto_in_a_bits_opcode; 
  assign a_io_enq_bits_size = auto_in_a_bits_size; 
  assign a_io_enq_bits_source = auto_in_a_bits_source; 
  assign a_io_deq_ready = _T_47 | _T_48; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  idle = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_15 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_117 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_161_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_33 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      idle <= 1'h1;
    end else begin
      if (_T_95) begin
        idle <= 1'h0;
      end
    end
    if (reset) begin
      _T_15 <= 4'h0;
    end else begin
      if (_T_6) begin
        if (_T_18) begin
          if (_T_13) begin
            _T_15 <= _T_11;
          end else begin
            _T_15 <= 4'h0;
          end
        end else begin
          _T_15 <= _T_17;
        end
      end
    end
    if (reset) begin
      _T_117 <= 4'h0;
    end else begin
      if (_T_119) begin
        if (_T_132) begin
          if (_T_31) begin
            _T_117 <= _T_30;
          end else begin
            _T_117 <= 4'h0;
          end
        end else begin
          _T_117 <= 4'h0;
        end
      end else begin
        _T_117 <= _T_158;
      end
    end
    if (reset) begin
      _T_161_1 <= 1'h0;
    end else begin
      if (_T_118) begin
        _T_161_1 <= _T_132;
      end
    end
    if (reset) begin
      _T_33 <= 4'h0;
    end else begin
      if (_T_25) begin
        if (da_first) begin
          if (_T_31) begin
            _T_33 <= _T_30;
          end else begin
            _T_33 <= 4'h0;
          end
        end else begin
          _T_33 <= _T_35;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_45) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Error.scala:28 assert (idle || da_first) // we only send Grant, never GrantData => simplified flow control below\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_45) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_152) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:70 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_152) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLFIFOFixer_1( 
  input         clock, 
  input         reset, 
  output        auto_in_a_ready, 
  input         auto_in_a_valid, 
  input  [2:0]  auto_in_a_bits_opcode, 
  input  [2:0]  auto_in_a_bits_param, 
  input  [3:0]  auto_in_a_bits_size, 
  input  [6:0]  auto_in_a_bits_source, 
  input  [31:0] auto_in_a_bits_address, 
  input  [7:0]  auto_in_a_bits_mask, 
  input  [63:0] auto_in_a_bits_data, 
  output        auto_in_c_ready, 
  input         auto_in_c_valid, 
  input  [2:0]  auto_in_c_bits_opcode, 
  input  [2:0]  auto_in_c_bits_param, 
  input  [3:0]  auto_in_c_bits_size, 
  input  [6:0]  auto_in_c_bits_source, 
  input  [31:0] auto_in_c_bits_address, 
  input         auto_in_c_bits_corrupt, 
  input         auto_in_d_ready, 
  output        auto_in_d_valid, 
  output [2:0]  auto_in_d_bits_opcode, 
  output [1:0]  auto_in_d_bits_param, 
  output [3:0]  auto_in_d_bits_size, 
  output [6:0]  auto_in_d_bits_source, 
  output        auto_in_d_bits_sink, 
  output        auto_in_d_bits_denied, 
  output [63:0] auto_in_d_bits_data, 
  output        auto_in_d_bits_corrupt, 
  output        auto_in_e_ready, 
  input         auto_in_e_valid, 
  input         auto_in_e_bits_sink, 
  input         auto_out_a_ready, 
  output        auto_out_a_valid, 
  output [2:0]  auto_out_a_bits_opcode, 
  output [2:0]  auto_out_a_bits_param, 
  output [3:0]  auto_out_a_bits_size, 
  output [6:0]  auto_out_a_bits_source, 
  output [31:0] auto_out_a_bits_address, 
  output [7:0]  auto_out_a_bits_mask, 
  output [63:0] auto_out_a_bits_data, 
  input         auto_out_c_ready, 
  output        auto_out_c_valid, 
  output [2:0]  auto_out_c_bits_opcode, 
  output [2:0]  auto_out_c_bits_param, 
  output [3:0]  auto_out_c_bits_size, 
  output [6:0]  auto_out_c_bits_source, 
  output [31:0] auto_out_c_bits_address, 
  output        auto_out_c_bits_corrupt, 
  output        auto_out_d_ready, 
  input         auto_out_d_valid, 
  input  [2:0]  auto_out_d_bits_opcode, 
  input  [1:0]  auto_out_d_bits_param, 
  input  [3:0]  auto_out_d_bits_size, 
  input  [6:0]  auto_out_d_bits_source, 
  input         auto_out_d_bits_sink, 
  input         auto_out_d_bits_denied, 
  input  [63:0] auto_out_d_bits_data, 
  input         auto_out_d_bits_corrupt, 
  input         auto_out_e_ready, 
  output        auto_out_e_valid, 
  output        auto_out_e_bits_sink 
);
  wire  TLMonitor_clock; 
  wire  TLMonitor_reset; 
  wire  TLMonitor_io_in_a_ready; 
  wire  TLMonitor_io_in_a_valid; 
  wire [2:0] TLMonitor_io_in_a_bits_opcode; 
  wire [2:0] TLMonitor_io_in_a_bits_param; 
  wire [3:0] TLMonitor_io_in_a_bits_size; 
  wire [6:0] TLMonitor_io_in_a_bits_source; 
  wire [31:0] TLMonitor_io_in_a_bits_address; 
  wire [7:0] TLMonitor_io_in_a_bits_mask; 
  wire  TLMonitor_io_in_c_ready; 
  wire  TLMonitor_io_in_c_valid; 
  wire [2:0] TLMonitor_io_in_c_bits_opcode; 
  wire [2:0] TLMonitor_io_in_c_bits_param; 
  wire [3:0] TLMonitor_io_in_c_bits_size; 
  wire [6:0] TLMonitor_io_in_c_bits_source; 
  wire [31:0] TLMonitor_io_in_c_bits_address; 
  wire  TLMonitor_io_in_c_bits_corrupt; 
  wire  TLMonitor_io_in_d_ready; 
  wire  TLMonitor_io_in_d_valid; 
  wire [2:0] TLMonitor_io_in_d_bits_opcode; 
  wire [1:0] TLMonitor_io_in_d_bits_param; 
  wire [3:0] TLMonitor_io_in_d_bits_size; 
  wire [6:0] TLMonitor_io_in_d_bits_source; 
  wire  TLMonitor_io_in_d_bits_sink; 
  wire  TLMonitor_io_in_d_bits_denied; 
  wire  TLMonitor_io_in_d_bits_corrupt; 
  wire  TLMonitor_io_in_e_ready; 
  wire  TLMonitor_io_in_e_valid; 
  wire  TLMonitor_io_in_e_bits_sink; 
  wire [32:0] _T_9; 
  wire [31:0] _T_13; 
  wire [32:0] _T_14; 
  wire [32:0] _T_15; 
  wire [32:0] _T_16; 
  wire  _T_17; 
  wire [31:0] _T_18; 
  wire [32:0] _T_19; 
  wire [32:0] _T_20; 
  wire [32:0] _T_21; 
  wire  _T_22; 
  wire [32:0] _T_25; 
  wire [32:0] _T_26; 
  wire  _T_27; 
  wire [1:0] _T_29; 
  wire [1:0] _T_30; 
  wire [1:0] _GEN_523; 
  wire [1:0] _T_31; 
  wire [1:0] _T_32; 
  wire  _T_34; 
  wire [2:0] _T_85; 
  wire  _T_86; 
  reg [4:0] _T_44; 
  reg [31:0] _RAND_0;
  wire  _T_47; 
  wire  _T_96; 
  reg  _T_77_16; 
  reg [31:0] _RAND_1;
  reg  _T_77_17; 
  reg [31:0] _RAND_2;
  wire  _T_97; 
  reg  _T_77_18; 
  reg [31:0] _RAND_3;
  wire  _T_98; 
  reg  _T_77_19; 
  reg [31:0] _RAND_4;
  wire  _T_99; 
  reg  _T_77_20; 
  reg [31:0] _RAND_5;
  wire  _T_100; 
  reg  _T_77_21; 
  reg [31:0] _RAND_6;
  wire  _T_101; 
  reg  _T_77_22; 
  reg [31:0] _RAND_7;
  wire  _T_102; 
  reg  _T_77_23; 
  reg [31:0] _RAND_8;
  wire  _T_103; 
  reg  _T_77_24; 
  reg [31:0] _RAND_9;
  wire  _T_104; 
  reg  _T_77_25; 
  reg [31:0] _RAND_10;
  wire  _T_105; 
  reg  _T_77_26; 
  reg [31:0] _RAND_11;
  wire  _T_106; 
  reg  _T_77_27; 
  reg [31:0] _RAND_12;
  wire  _T_107; 
  reg  _T_77_28; 
  reg [31:0] _RAND_13;
  wire  _T_108; 
  reg  _T_77_29; 
  reg [31:0] _RAND_14;
  wire  _T_109; 
  reg  _T_77_30; 
  reg [31:0] _RAND_15;
  wire  _T_110; 
  reg  _T_77_31; 
  reg [31:0] _RAND_16;
  wire  _T_111; 
  wire  _T_112; 
  reg [1:0] _T_95; 
  reg [31:0] _RAND_17;
  wire  _T_113; 
  wire  _T_114; 
  wire  _T_115; 
  wire  _T_119; 
  wire  _T_129; 
  reg  _T_77_32; 
  reg [31:0] _RAND_18;
  reg  _T_77_33; 
  reg [31:0] _RAND_19;
  wire  _T_130; 
  reg  _T_77_34; 
  reg [31:0] _RAND_20;
  wire  _T_131; 
  reg  _T_77_35; 
  reg [31:0] _RAND_21;
  wire  _T_132; 
  reg  _T_77_36; 
  reg [31:0] _RAND_22;
  wire  _T_133; 
  reg  _T_77_37; 
  reg [31:0] _RAND_23;
  wire  _T_134; 
  reg  _T_77_38; 
  reg [31:0] _RAND_24;
  wire  _T_135; 
  reg  _T_77_39; 
  reg [31:0] _RAND_25;
  wire  _T_136; 
  reg  _T_77_40; 
  reg [31:0] _RAND_26;
  wire  _T_137; 
  reg  _T_77_41; 
  reg [31:0] _RAND_27;
  wire  _T_138; 
  reg  _T_77_42; 
  reg [31:0] _RAND_28;
  wire  _T_139; 
  reg  _T_77_43; 
  reg [31:0] _RAND_29;
  wire  _T_140; 
  reg  _T_77_44; 
  reg [31:0] _RAND_30;
  wire  _T_141; 
  reg  _T_77_45; 
  reg [31:0] _RAND_31;
  wire  _T_142; 
  reg  _T_77_46; 
  reg [31:0] _RAND_32;
  wire  _T_143; 
  reg  _T_77_47; 
  reg [31:0] _RAND_33;
  wire  _T_144; 
  wire  _T_145; 
  reg [1:0] _T_128; 
  reg [31:0] _RAND_34;
  wire  _T_146; 
  wire  _T_147; 
  wire  _T_148; 
  wire  _T_315; 
  wire  _T_152; 
  wire  _T_162; 
  reg  _T_77_48; 
  reg [31:0] _RAND_35;
  reg  _T_77_49; 
  reg [31:0] _RAND_36;
  wire  _T_163; 
  reg  _T_77_50; 
  reg [31:0] _RAND_37;
  wire  _T_164; 
  reg  _T_77_51; 
  reg [31:0] _RAND_38;
  wire  _T_165; 
  reg  _T_77_52; 
  reg [31:0] _RAND_39;
  wire  _T_166; 
  reg  _T_77_53; 
  reg [31:0] _RAND_40;
  wire  _T_167; 
  reg  _T_77_54; 
  reg [31:0] _RAND_41;
  wire  _T_168; 
  reg  _T_77_55; 
  reg [31:0] _RAND_42;
  wire  _T_169; 
  reg  _T_77_56; 
  reg [31:0] _RAND_43;
  wire  _T_170; 
  reg  _T_77_57; 
  reg [31:0] _RAND_44;
  wire  _T_171; 
  reg  _T_77_58; 
  reg [31:0] _RAND_45;
  wire  _T_172; 
  reg  _T_77_59; 
  reg [31:0] _RAND_46;
  wire  _T_173; 
  reg  _T_77_60; 
  reg [31:0] _RAND_47;
  wire  _T_174; 
  reg  _T_77_61; 
  reg [31:0] _RAND_48;
  wire  _T_175; 
  reg  _T_77_62; 
  reg [31:0] _RAND_49;
  wire  _T_176; 
  reg  _T_77_63; 
  reg [31:0] _RAND_50;
  wire  _T_177; 
  wire  _T_178; 
  reg [1:0] _T_161; 
  reg [31:0] _RAND_51;
  wire  _T_179; 
  wire  _T_180; 
  wire  _T_181; 
  wire  _T_316; 
  wire  _T_185; 
  wire  _T_195; 
  reg  _T_77_64; 
  reg [31:0] _RAND_52;
  reg  _T_77_65; 
  reg [31:0] _RAND_53;
  wire  _T_196; 
  reg  _T_77_66; 
  reg [31:0] _RAND_54;
  wire  _T_197; 
  reg  _T_77_67; 
  reg [31:0] _RAND_55;
  wire  _T_198; 
  reg  _T_77_68; 
  reg [31:0] _RAND_56;
  wire  _T_199; 
  reg  _T_77_69; 
  reg [31:0] _RAND_57;
  wire  _T_200; 
  reg  _T_77_70; 
  reg [31:0] _RAND_58;
  wire  _T_201; 
  reg  _T_77_71; 
  reg [31:0] _RAND_59;
  wire  _T_202; 
  reg  _T_77_72; 
  reg [31:0] _RAND_60;
  wire  _T_203; 
  reg  _T_77_73; 
  reg [31:0] _RAND_61;
  wire  _T_204; 
  reg  _T_77_74; 
  reg [31:0] _RAND_62;
  wire  _T_205; 
  reg  _T_77_75; 
  reg [31:0] _RAND_63;
  wire  _T_206; 
  reg  _T_77_76; 
  reg [31:0] _RAND_64;
  wire  _T_207; 
  reg  _T_77_77; 
  reg [31:0] _RAND_65;
  wire  _T_208; 
  reg  _T_77_78; 
  reg [31:0] _RAND_66;
  wire  _T_209; 
  reg  _T_77_79; 
  reg [31:0] _RAND_67;
  wire  _T_210; 
  wire  _T_211; 
  reg [1:0] _T_194; 
  reg [31:0] _RAND_68;
  wire  _T_212; 
  wire  _T_213; 
  wire  _T_214; 
  wire  _T_317; 
  wire  _T_218; 
  wire  _T_228; 
  reg  _T_77_80; 
  reg [31:0] _RAND_69;
  reg  _T_77_81; 
  reg [31:0] _RAND_70;
  wire  _T_229; 
  reg  _T_77_82; 
  reg [31:0] _RAND_71;
  wire  _T_230; 
  reg  _T_77_83; 
  reg [31:0] _RAND_72;
  wire  _T_231; 
  reg  _T_77_84; 
  reg [31:0] _RAND_73;
  wire  _T_232; 
  reg  _T_77_85; 
  reg [31:0] _RAND_74;
  wire  _T_233; 
  reg  _T_77_86; 
  reg [31:0] _RAND_75;
  wire  _T_234; 
  reg  _T_77_87; 
  reg [31:0] _RAND_76;
  wire  _T_235; 
  reg  _T_77_88; 
  reg [31:0] _RAND_77;
  wire  _T_236; 
  reg  _T_77_89; 
  reg [31:0] _RAND_78;
  wire  _T_237; 
  reg  _T_77_90; 
  reg [31:0] _RAND_79;
  wire  _T_238; 
  reg  _T_77_91; 
  reg [31:0] _RAND_80;
  wire  _T_239; 
  reg  _T_77_92; 
  reg [31:0] _RAND_81;
  wire  _T_240; 
  reg  _T_77_93; 
  reg [31:0] _RAND_82;
  wire  _T_241; 
  reg  _T_77_94; 
  reg [31:0] _RAND_83;
  wire  _T_242; 
  reg  _T_77_95; 
  reg [31:0] _RAND_84;
  wire  _T_243; 
  wire  _T_244; 
  reg [1:0] _T_227; 
  reg [31:0] _RAND_85;
  wire  _T_245; 
  wire  _T_246; 
  wire  _T_247; 
  wire  _T_318; 
  wire  _T_251; 
  wire  _T_261; 
  reg  _T_77_96; 
  reg [31:0] _RAND_86;
  reg  _T_77_97; 
  reg [31:0] _RAND_87;
  wire  _T_262; 
  reg  _T_77_98; 
  reg [31:0] _RAND_88;
  wire  _T_263; 
  reg  _T_77_99; 
  reg [31:0] _RAND_89;
  wire  _T_264; 
  reg  _T_77_100; 
  reg [31:0] _RAND_90;
  wire  _T_265; 
  reg  _T_77_101; 
  reg [31:0] _RAND_91;
  wire  _T_266; 
  reg  _T_77_102; 
  reg [31:0] _RAND_92;
  wire  _T_267; 
  reg  _T_77_103; 
  reg [31:0] _RAND_93;
  wire  _T_268; 
  reg  _T_77_104; 
  reg [31:0] _RAND_94;
  wire  _T_269; 
  reg  _T_77_105; 
  reg [31:0] _RAND_95;
  wire  _T_270; 
  reg  _T_77_106; 
  reg [31:0] _RAND_96;
  wire  _T_271; 
  reg  _T_77_107; 
  reg [31:0] _RAND_97;
  wire  _T_272; 
  reg  _T_77_108; 
  reg [31:0] _RAND_98;
  wire  _T_273; 
  reg  _T_77_109; 
  reg [31:0] _RAND_99;
  wire  _T_274; 
  reg  _T_77_110; 
  reg [31:0] _RAND_100;
  wire  _T_275; 
  reg  _T_77_111; 
  reg [31:0] _RAND_101;
  wire  _T_276; 
  wire  _T_277; 
  reg [1:0] _T_260; 
  reg [31:0] _RAND_102;
  wire  _T_278; 
  wire  _T_279; 
  wire  _T_280; 
  wire  _T_319; 
  wire  _T_284; 
  wire  _T_294; 
  reg  _T_77_112; 
  reg [31:0] _RAND_103;
  reg  _T_77_113; 
  reg [31:0] _RAND_104;
  wire  _T_295; 
  reg  _T_77_114; 
  reg [31:0] _RAND_105;
  wire  _T_296; 
  reg  _T_77_115; 
  reg [31:0] _RAND_106;
  wire  _T_297; 
  reg  _T_77_116; 
  reg [31:0] _RAND_107;
  wire  _T_298; 
  reg  _T_77_117; 
  reg [31:0] _RAND_108;
  wire  _T_299; 
  reg  _T_77_118; 
  reg [31:0] _RAND_109;
  wire  _T_300; 
  reg  _T_77_119; 
  reg [31:0] _RAND_110;
  wire  _T_301; 
  reg  _T_77_120; 
  reg [31:0] _RAND_111;
  wire  _T_302; 
  reg  _T_77_121; 
  reg [31:0] _RAND_112;
  wire  _T_303; 
  reg  _T_77_122; 
  reg [31:0] _RAND_113;
  wire  _T_304; 
  reg  _T_77_123; 
  reg [31:0] _RAND_114;
  wire  _T_305; 
  reg  _T_77_124; 
  reg [31:0] _RAND_115;
  wire  _T_306; 
  reg  _T_77_125; 
  reg [31:0] _RAND_116;
  wire  _T_307; 
  reg  _T_77_126; 
  reg [31:0] _RAND_117;
  wire  _T_308; 
  reg  _T_77_127; 
  reg [31:0] _RAND_118;
  wire  _T_309; 
  wire  _T_310; 
  reg [1:0] _T_293; 
  reg [31:0] _RAND_119;
  wire  _T_311; 
  wire  _T_312; 
  wire  _T_313; 
  wire  _T_320; 
  wire  _T_324; 
  wire  _T_326; 
  wire  _T_35; 
  wire [22:0] _T_37; 
  wire [7:0] _T_38; 
  wire [7:0] _T_39; 
  wire [4:0] _T_40; 
  wire  _T_41; 
  wire  _T_42; 
  wire [4:0] _T_46; 
  wire  _T_55; 
  wire [22:0] _T_57; 
  wire [7:0] _T_58; 
  wire [7:0] _T_59; 
  wire [4:0] _T_60; 
  wire  _T_61; 
  reg [4:0] _T_63; 
  reg [31:0] _RAND_120;
  wire [4:0] _T_65; 
  wire  _T_66; 
  wire  _T_74; 
  wire  _T_75; 
  wire  _T_79; 
  wire  _T_82; 
  wire  _T_92; 
  wire  _T_125; 
  wire  _T_158; 
  wire  _T_191; 
  wire  _T_224; 
  wire  _T_257; 
  wire  _T_290; 
  dual_TLMonitor_15 dual_TLMonitor ( 
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_c_ready(TLMonitor_io_in_c_ready),
    .io_in_c_valid(TLMonitor_io_in_c_valid),
    .io_in_c_bits_opcode(TLMonitor_io_in_c_bits_opcode),
    .io_in_c_bits_param(TLMonitor_io_in_c_bits_param),
    .io_in_c_bits_size(TLMonitor_io_in_c_bits_size),
    .io_in_c_bits_source(TLMonitor_io_in_c_bits_source),
    .io_in_c_bits_address(TLMonitor_io_in_c_bits_address),
    .io_in_c_bits_corrupt(TLMonitor_io_in_c_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt),
    .io_in_e_ready(TLMonitor_io_in_e_ready),
    .io_in_e_valid(TLMonitor_io_in_e_valid),
    .io_in_e_bits_sink(TLMonitor_io_in_e_bits_sink)
  );
  assign _T_9 = {1'b0,$signed(auto_in_a_bits_address)}; 
  assign _T_13 = auto_in_a_bits_address ^ 32'h80000000; 
  assign _T_14 = {1'b0,$signed(_T_13)}; 
  assign _T_15 = $signed(_T_14) & $signed(33'sh80000000); 
  assign _T_16 = $signed(_T_15); 
  assign _T_17 = $signed(_T_16) == $signed(33'sh0); 
  assign _T_18 = auto_in_a_bits_address ^ 32'h40000000; 
  assign _T_19 = {1'b0,$signed(_T_18)}; 
  assign _T_20 = $signed(_T_19) & $signed(33'shc0000000); 
  assign _T_21 = $signed(_T_20); 
  assign _T_22 = $signed(_T_21) == $signed(33'sh0); 
  assign _T_25 = $signed(_T_9) & $signed(33'shc0000000); 
  assign _T_26 = $signed(_T_25); 
  assign _T_27 = $signed(_T_26) == $signed(33'sh0); 
  assign _T_29 = _T_22 ? 2'h2 : 2'h0; 
  assign _T_30 = _T_27 ? 2'h3 : 2'h0; 
  assign _GEN_523 = {{1'd0}, _T_17}; 
  assign _T_31 = _GEN_523 | _T_29; 
  assign _T_32 = _T_31 | _T_30; 
  assign _T_34 = _T_32 == 2'h0; 
  assign _T_85 = auto_in_a_bits_source[6:4]; 
  assign _T_86 = _T_85 == 3'h1; 
  assign _T_47 = _T_44 == 5'h0; 
  assign _T_96 = _T_86 & _T_47; 
  assign _T_97 = _T_77_16 | _T_77_17; 
  assign _T_98 = _T_97 | _T_77_18; 
  assign _T_99 = _T_98 | _T_77_19; 
  assign _T_100 = _T_99 | _T_77_20; 
  assign _T_101 = _T_100 | _T_77_21; 
  assign _T_102 = _T_101 | _T_77_22; 
  assign _T_103 = _T_102 | _T_77_23; 
  assign _T_104 = _T_103 | _T_77_24; 
  assign _T_105 = _T_104 | _T_77_25; 
  assign _T_106 = _T_105 | _T_77_26; 
  assign _T_107 = _T_106 | _T_77_27; 
  assign _T_108 = _T_107 | _T_77_28; 
  assign _T_109 = _T_108 | _T_77_29; 
  assign _T_110 = _T_109 | _T_77_30; 
  assign _T_111 = _T_110 | _T_77_31; 
  assign _T_112 = _T_96 & _T_111; 
  assign _T_113 = _T_95 != _T_32; 
  assign _T_114 = _T_34 | _T_113; 
  assign _T_115 = _T_112 & _T_114; 
  assign _T_119 = _T_85 == 3'h2; 
  assign _T_129 = _T_119 & _T_47; 
  assign _T_130 = _T_77_32 | _T_77_33; 
  assign _T_131 = _T_130 | _T_77_34; 
  assign _T_132 = _T_131 | _T_77_35; 
  assign _T_133 = _T_132 | _T_77_36; 
  assign _T_134 = _T_133 | _T_77_37; 
  assign _T_135 = _T_134 | _T_77_38; 
  assign _T_136 = _T_135 | _T_77_39; 
  assign _T_137 = _T_136 | _T_77_40; 
  assign _T_138 = _T_137 | _T_77_41; 
  assign _T_139 = _T_138 | _T_77_42; 
  assign _T_140 = _T_139 | _T_77_43; 
  assign _T_141 = _T_140 | _T_77_44; 
  assign _T_142 = _T_141 | _T_77_45; 
  assign _T_143 = _T_142 | _T_77_46; 
  assign _T_144 = _T_143 | _T_77_47; 
  assign _T_145 = _T_129 & _T_144; 
  assign _T_146 = _T_128 != _T_32; 
  assign _T_147 = _T_34 | _T_146; 
  assign _T_148 = _T_145 & _T_147; 
  assign _T_315 = _T_115 | _T_148; 
  assign _T_152 = _T_85 == 3'h3; 
  assign _T_162 = _T_152 & _T_47; 
  assign _T_163 = _T_77_48 | _T_77_49; 
  assign _T_164 = _T_163 | _T_77_50; 
  assign _T_165 = _T_164 | _T_77_51; 
  assign _T_166 = _T_165 | _T_77_52; 
  assign _T_167 = _T_166 | _T_77_53; 
  assign _T_168 = _T_167 | _T_77_54; 
  assign _T_169 = _T_168 | _T_77_55; 
  assign _T_170 = _T_169 | _T_77_56; 
  assign _T_171 = _T_170 | _T_77_57; 
  assign _T_172 = _T_171 | _T_77_58; 
  assign _T_173 = _T_172 | _T_77_59; 
  assign _T_174 = _T_173 | _T_77_60; 
  assign _T_175 = _T_174 | _T_77_61; 
  assign _T_176 = _T_175 | _T_77_62; 
  assign _T_177 = _T_176 | _T_77_63; 
  assign _T_178 = _T_162 & _T_177; 
  assign _T_179 = _T_161 != _T_32; 
  assign _T_180 = _T_34 | _T_179; 
  assign _T_181 = _T_178 & _T_180; 
  assign _T_316 = _T_315 | _T_181; 
  assign _T_185 = _T_85 == 3'h4; 
  assign _T_195 = _T_185 & _T_47; 
  assign _T_196 = _T_77_64 | _T_77_65; 
  assign _T_197 = _T_196 | _T_77_66; 
  assign _T_198 = _T_197 | _T_77_67; 
  assign _T_199 = _T_198 | _T_77_68; 
  assign _T_200 = _T_199 | _T_77_69; 
  assign _T_201 = _T_200 | _T_77_70; 
  assign _T_202 = _T_201 | _T_77_71; 
  assign _T_203 = _T_202 | _T_77_72; 
  assign _T_204 = _T_203 | _T_77_73; 
  assign _T_205 = _T_204 | _T_77_74; 
  assign _T_206 = _T_205 | _T_77_75; 
  assign _T_207 = _T_206 | _T_77_76; 
  assign _T_208 = _T_207 | _T_77_77; 
  assign _T_209 = _T_208 | _T_77_78; 
  assign _T_210 = _T_209 | _T_77_79; 
  assign _T_211 = _T_195 & _T_210; 
  assign _T_212 = _T_194 != _T_32; 
  assign _T_213 = _T_34 | _T_212; 
  assign _T_214 = _T_211 & _T_213; 
  assign _T_317 = _T_316 | _T_214; 
  assign _T_218 = _T_85 == 3'h5; 
  assign _T_228 = _T_218 & _T_47; 
  assign _T_229 = _T_77_80 | _T_77_81; 
  assign _T_230 = _T_229 | _T_77_82; 
  assign _T_231 = _T_230 | _T_77_83; 
  assign _T_232 = _T_231 | _T_77_84; 
  assign _T_233 = _T_232 | _T_77_85; 
  assign _T_234 = _T_233 | _T_77_86; 
  assign _T_235 = _T_234 | _T_77_87; 
  assign _T_236 = _T_235 | _T_77_88; 
  assign _T_237 = _T_236 | _T_77_89; 
  assign _T_238 = _T_237 | _T_77_90; 
  assign _T_239 = _T_238 | _T_77_91; 
  assign _T_240 = _T_239 | _T_77_92; 
  assign _T_241 = _T_240 | _T_77_93; 
  assign _T_242 = _T_241 | _T_77_94; 
  assign _T_243 = _T_242 | _T_77_95; 
  assign _T_244 = _T_228 & _T_243; 
  assign _T_245 = _T_227 != _T_32; 
  assign _T_246 = _T_34 | _T_245; 
  assign _T_247 = _T_244 & _T_246; 
  assign _T_318 = _T_317 | _T_247; 
  assign _T_251 = _T_85 == 3'h6; 
  assign _T_261 = _T_251 & _T_47; 
  assign _T_262 = _T_77_96 | _T_77_97; 
  assign _T_263 = _T_262 | _T_77_98; 
  assign _T_264 = _T_263 | _T_77_99; 
  assign _T_265 = _T_264 | _T_77_100; 
  assign _T_266 = _T_265 | _T_77_101; 
  assign _T_267 = _T_266 | _T_77_102; 
  assign _T_268 = _T_267 | _T_77_103; 
  assign _T_269 = _T_268 | _T_77_104; 
  assign _T_270 = _T_269 | _T_77_105; 
  assign _T_271 = _T_270 | _T_77_106; 
  assign _T_272 = _T_271 | _T_77_107; 
  assign _T_273 = _T_272 | _T_77_108; 
  assign _T_274 = _T_273 | _T_77_109; 
  assign _T_275 = _T_274 | _T_77_110; 
  assign _T_276 = _T_275 | _T_77_111; 
  assign _T_277 = _T_261 & _T_276; 
  assign _T_278 = _T_260 != _T_32; 
  assign _T_279 = _T_34 | _T_278; 
  assign _T_280 = _T_277 & _T_279; 
  assign _T_319 = _T_318 | _T_280; 
  assign _T_284 = _T_85 == 3'h7; 
  assign _T_294 = _T_284 & _T_47; 
  assign _T_295 = _T_77_112 | _T_77_113; 
  assign _T_296 = _T_295 | _T_77_114; 
  assign _T_297 = _T_296 | _T_77_115; 
  assign _T_298 = _T_297 | _T_77_116; 
  assign _T_299 = _T_298 | _T_77_117; 
  assign _T_300 = _T_299 | _T_77_118; 
  assign _T_301 = _T_300 | _T_77_119; 
  assign _T_302 = _T_301 | _T_77_120; 
  assign _T_303 = _T_302 | _T_77_121; 
  assign _T_304 = _T_303 | _T_77_122; 
  assign _T_305 = _T_304 | _T_77_123; 
  assign _T_306 = _T_305 | _T_77_124; 
  assign _T_307 = _T_306 | _T_77_125; 
  assign _T_308 = _T_307 | _T_77_126; 
  assign _T_309 = _T_308 | _T_77_127; 
  assign _T_310 = _T_294 & _T_309; 
  assign _T_311 = _T_293 != _T_32; 
  assign _T_312 = _T_34 | _T_311; 
  assign _T_313 = _T_310 & _T_312; 
  assign _T_320 = _T_319 | _T_313; 
  assign _T_324 = _T_320 == 1'h0; 
  assign _T_326 = auto_out_a_ready & _T_324; 
  assign _T_35 = _T_326 & auto_in_a_valid; 
  assign _T_37 = 23'hff << auto_in_a_bits_size; 
  assign _T_38 = _T_37[7:0]; 
  assign _T_39 = ~ _T_38; 
  assign _T_40 = _T_39[7:3]; 
  assign _T_41 = auto_in_a_bits_opcode[2]; 
  assign _T_42 = _T_41 == 1'h0; 
  assign _T_46 = _T_44 - 5'h1; 
  assign _T_55 = auto_in_d_ready & auto_out_d_valid; 
  assign _T_57 = 23'hff << auto_out_d_bits_size; 
  assign _T_58 = _T_57[7:0]; 
  assign _T_59 = ~ _T_58; 
  assign _T_60 = _T_59[7:3]; 
  assign _T_61 = auto_out_d_bits_opcode[0]; 
  assign _T_65 = _T_63 - 5'h1; 
  assign _T_66 = _T_63 == 5'h0; 
  assign _T_74 = auto_out_d_bits_opcode != 3'h6; 
  assign _T_75 = _T_66 & _T_74; 
  assign _T_79 = _T_47 & _T_35; 
  assign _T_82 = _T_75 & _T_55; 
  assign _T_92 = _T_35 & _T_86; 
  assign _T_125 = _T_35 & _T_119; 
  assign _T_158 = _T_35 & _T_152; 
  assign _T_191 = _T_35 & _T_185; 
  assign _T_224 = _T_35 & _T_218; 
  assign _T_257 = _T_35 & _T_251; 
  assign _T_290 = _T_35 & _T_284; 
  assign auto_in_a_ready = auto_out_a_ready & _T_324; 
  assign auto_in_c_ready = auto_out_c_ready; 
  assign auto_in_d_valid = auto_out_d_valid; 
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; 
  assign auto_in_d_bits_param = auto_out_d_bits_param; 
  assign auto_in_d_bits_size = auto_out_d_bits_size; 
  assign auto_in_d_bits_source = auto_out_d_bits_source; 
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; 
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; 
  assign auto_in_d_bits_data = auto_out_d_bits_data; 
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; 
  assign auto_in_e_ready = auto_out_e_ready; 
  assign auto_out_a_valid = auto_in_a_valid & _T_324; 
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; 
  assign auto_out_a_bits_param = auto_in_a_bits_param; 
  assign auto_out_a_bits_size = auto_in_a_bits_size; 
  assign auto_out_a_bits_source = auto_in_a_bits_source; 
  assign auto_out_a_bits_address = auto_in_a_bits_address; 
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; 
  assign auto_out_a_bits_data = auto_in_a_bits_data; 
  assign auto_out_c_valid = auto_in_c_valid; 
  assign auto_out_c_bits_opcode = auto_in_c_bits_opcode; 
  assign auto_out_c_bits_param = auto_in_c_bits_param; 
  assign auto_out_c_bits_size = auto_in_c_bits_size; 
  assign auto_out_c_bits_source = auto_in_c_bits_source; 
  assign auto_out_c_bits_address = auto_in_c_bits_address; 
  assign auto_out_c_bits_corrupt = auto_in_c_bits_corrupt; 
  assign auto_out_d_ready = auto_in_d_ready; 
  assign auto_out_e_valid = auto_in_e_valid; 
  assign auto_out_e_bits_sink = auto_in_e_bits_sink; 
  assign TLMonitor_clock = clock; 
  assign TLMonitor_reset = reset; 
  assign TLMonitor_io_in_a_ready = auto_out_a_ready & _T_324; 
  assign TLMonitor_io_in_a_valid = auto_in_a_valid; 
  assign TLMonitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; 
  assign TLMonitor_io_in_a_bits_param = auto_in_a_bits_param; 
  assign TLMonitor_io_in_a_bits_size = auto_in_a_bits_size; 
  assign TLMonitor_io_in_a_bits_source = auto_in_a_bits_source; 
  assign TLMonitor_io_in_a_bits_address = auto_in_a_bits_address; 
  assign TLMonitor_io_in_a_bits_mask = auto_in_a_bits_mask; 
  assign TLMonitor_io_in_c_ready = auto_out_c_ready; 
  assign TLMonitor_io_in_c_valid = auto_in_c_valid; 
  assign TLMonitor_io_in_c_bits_opcode = auto_in_c_bits_opcode; 
  assign TLMonitor_io_in_c_bits_param = auto_in_c_bits_param; 
  assign TLMonitor_io_in_c_bits_size = auto_in_c_bits_size; 
  assign TLMonitor_io_in_c_bits_source = auto_in_c_bits_source; 
  assign TLMonitor_io_in_c_bits_address = auto_in_c_bits_address; 
  assign TLMonitor_io_in_c_bits_corrupt = auto_in_c_bits_corrupt; 
  assign TLMonitor_io_in_d_ready = auto_in_d_ready; 
  assign TLMonitor_io_in_d_valid = auto_out_d_valid; 
  assign TLMonitor_io_in_d_bits_opcode = auto_out_d_bits_opcode; 
  assign TLMonitor_io_in_d_bits_param = auto_out_d_bits_param; 
  assign TLMonitor_io_in_d_bits_size = auto_out_d_bits_size; 
  assign TLMonitor_io_in_d_bits_source = auto_out_d_bits_source; 
  assign TLMonitor_io_in_d_bits_sink = auto_out_d_bits_sink; 
  assign TLMonitor_io_in_d_bits_denied = auto_out_d_bits_denied; 
  assign TLMonitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; 
  assign TLMonitor_io_in_e_ready = auto_out_e_ready; 
  assign TLMonitor_io_in_e_valid = auto_in_e_valid; 
  assign TLMonitor_io_in_e_bits_sink = auto_in_e_bits_sink; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_44 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_77_16 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_77_17 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_77_18 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_77_19 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_77_20 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_77_21 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_77_22 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_77_23 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_77_24 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_77_25 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_77_26 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_77_27 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_77_28 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_77_29 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_77_30 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_77_31 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_95 = _RAND_17[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_77_32 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_77_33 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_77_34 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_77_35 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_77_36 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_77_37 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_77_38 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_77_39 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_77_40 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_77_41 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_77_42 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_77_43 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_77_44 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_77_45 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_77_46 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_77_47 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_128 = _RAND_34[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_77_48 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_77_49 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_77_50 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_77_51 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_77_52 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_77_53 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_77_54 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_77_55 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_77_56 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_77_57 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_77_58 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_77_59 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_77_60 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_77_61 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_77_62 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_77_63 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_161 = _RAND_51[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_77_64 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_77_65 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_77_66 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_77_67 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_77_68 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_77_69 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_77_70 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_77_71 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_77_72 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_77_73 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_77_74 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_77_75 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_77_76 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_77_77 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_77_78 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_77_79 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_194 = _RAND_68[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_77_80 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_77_81 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_77_82 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_77_83 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_77_84 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_77_85 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_77_86 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_77_87 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_77_88 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_77_89 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_77_90 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_77_91 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_77_92 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_77_93 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_77_94 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_77_95 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_227 = _RAND_85[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_77_96 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_77_97 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_77_98 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_77_99 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_77_100 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_77_101 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_77_102 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_77_103 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_77_104 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_77_105 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_77_106 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_77_107 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_77_108 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_77_109 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_77_110 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_77_111 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_260 = _RAND_102[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_77_112 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_77_113 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_77_114 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_77_115 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_77_116 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_77_117 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_77_118 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_77_119 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_77_120 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_77_121 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_77_122 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_77_123 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_77_124 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_77_125 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_77_126 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_77_127 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_293 = _RAND_119[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_63 = _RAND_120[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_44 <= 5'h0;
    end else begin
      if (_T_35) begin
        if (_T_47) begin
          if (_T_42) begin
            _T_44 <= _T_40;
          end else begin
            _T_44 <= 5'h0;
          end
        end else begin
          _T_44 <= _T_46;
        end
      end
    end
    if (reset) begin
      _T_77_16 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h10 == auto_out_d_bits_source) begin
          _T_77_16 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h10 == auto_in_a_bits_source) begin
              _T_77_16 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h10 == auto_in_a_bits_source) begin
            _T_77_16 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_17 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h11 == auto_out_d_bits_source) begin
          _T_77_17 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h11 == auto_in_a_bits_source) begin
              _T_77_17 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h11 == auto_in_a_bits_source) begin
            _T_77_17 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_18 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h12 == auto_out_d_bits_source) begin
          _T_77_18 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h12 == auto_in_a_bits_source) begin
              _T_77_18 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h12 == auto_in_a_bits_source) begin
            _T_77_18 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_19 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h13 == auto_out_d_bits_source) begin
          _T_77_19 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h13 == auto_in_a_bits_source) begin
              _T_77_19 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h13 == auto_in_a_bits_source) begin
            _T_77_19 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_20 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h14 == auto_out_d_bits_source) begin
          _T_77_20 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h14 == auto_in_a_bits_source) begin
              _T_77_20 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h14 == auto_in_a_bits_source) begin
            _T_77_20 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_21 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h15 == auto_out_d_bits_source) begin
          _T_77_21 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h15 == auto_in_a_bits_source) begin
              _T_77_21 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h15 == auto_in_a_bits_source) begin
            _T_77_21 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_22 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h16 == auto_out_d_bits_source) begin
          _T_77_22 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h16 == auto_in_a_bits_source) begin
              _T_77_22 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h16 == auto_in_a_bits_source) begin
            _T_77_22 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_23 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h17 == auto_out_d_bits_source) begin
          _T_77_23 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h17 == auto_in_a_bits_source) begin
              _T_77_23 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h17 == auto_in_a_bits_source) begin
            _T_77_23 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_24 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h18 == auto_out_d_bits_source) begin
          _T_77_24 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h18 == auto_in_a_bits_source) begin
              _T_77_24 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h18 == auto_in_a_bits_source) begin
            _T_77_24 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_25 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h19 == auto_out_d_bits_source) begin
          _T_77_25 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h19 == auto_in_a_bits_source) begin
              _T_77_25 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h19 == auto_in_a_bits_source) begin
            _T_77_25 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_26 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h1a == auto_out_d_bits_source) begin
          _T_77_26 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h1a == auto_in_a_bits_source) begin
              _T_77_26 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h1a == auto_in_a_bits_source) begin
            _T_77_26 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_27 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h1b == auto_out_d_bits_source) begin
          _T_77_27 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h1b == auto_in_a_bits_source) begin
              _T_77_27 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h1b == auto_in_a_bits_source) begin
            _T_77_27 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_28 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h1c == auto_out_d_bits_source) begin
          _T_77_28 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h1c == auto_in_a_bits_source) begin
              _T_77_28 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h1c == auto_in_a_bits_source) begin
            _T_77_28 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_29 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h1d == auto_out_d_bits_source) begin
          _T_77_29 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h1d == auto_in_a_bits_source) begin
              _T_77_29 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h1d == auto_in_a_bits_source) begin
            _T_77_29 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_30 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h1e == auto_out_d_bits_source) begin
          _T_77_30 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h1e == auto_in_a_bits_source) begin
              _T_77_30 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h1e == auto_in_a_bits_source) begin
            _T_77_30 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_31 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h1f == auto_out_d_bits_source) begin
          _T_77_31 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h1f == auto_in_a_bits_source) begin
              _T_77_31 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h1f == auto_in_a_bits_source) begin
            _T_77_31 <= 1'h1;
          end
        end
      end
    end
    if (_T_92) begin
      _T_95 <= _T_32;
    end
    if (reset) begin
      _T_77_32 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h20 == auto_out_d_bits_source) begin
          _T_77_32 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h20 == auto_in_a_bits_source) begin
              _T_77_32 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h20 == auto_in_a_bits_source) begin
            _T_77_32 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_33 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h21 == auto_out_d_bits_source) begin
          _T_77_33 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h21 == auto_in_a_bits_source) begin
              _T_77_33 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h21 == auto_in_a_bits_source) begin
            _T_77_33 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_34 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h22 == auto_out_d_bits_source) begin
          _T_77_34 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h22 == auto_in_a_bits_source) begin
              _T_77_34 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h22 == auto_in_a_bits_source) begin
            _T_77_34 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_35 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h23 == auto_out_d_bits_source) begin
          _T_77_35 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h23 == auto_in_a_bits_source) begin
              _T_77_35 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h23 == auto_in_a_bits_source) begin
            _T_77_35 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_36 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h24 == auto_out_d_bits_source) begin
          _T_77_36 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h24 == auto_in_a_bits_source) begin
              _T_77_36 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h24 == auto_in_a_bits_source) begin
            _T_77_36 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_37 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h25 == auto_out_d_bits_source) begin
          _T_77_37 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h25 == auto_in_a_bits_source) begin
              _T_77_37 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h25 == auto_in_a_bits_source) begin
            _T_77_37 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_38 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h26 == auto_out_d_bits_source) begin
          _T_77_38 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h26 == auto_in_a_bits_source) begin
              _T_77_38 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h26 == auto_in_a_bits_source) begin
            _T_77_38 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_39 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h27 == auto_out_d_bits_source) begin
          _T_77_39 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h27 == auto_in_a_bits_source) begin
              _T_77_39 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h27 == auto_in_a_bits_source) begin
            _T_77_39 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_40 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h28 == auto_out_d_bits_source) begin
          _T_77_40 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h28 == auto_in_a_bits_source) begin
              _T_77_40 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h28 == auto_in_a_bits_source) begin
            _T_77_40 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_41 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h29 == auto_out_d_bits_source) begin
          _T_77_41 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h29 == auto_in_a_bits_source) begin
              _T_77_41 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h29 == auto_in_a_bits_source) begin
            _T_77_41 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_42 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h2a == auto_out_d_bits_source) begin
          _T_77_42 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h2a == auto_in_a_bits_source) begin
              _T_77_42 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h2a == auto_in_a_bits_source) begin
            _T_77_42 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_43 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h2b == auto_out_d_bits_source) begin
          _T_77_43 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h2b == auto_in_a_bits_source) begin
              _T_77_43 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h2b == auto_in_a_bits_source) begin
            _T_77_43 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_44 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h2c == auto_out_d_bits_source) begin
          _T_77_44 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h2c == auto_in_a_bits_source) begin
              _T_77_44 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h2c == auto_in_a_bits_source) begin
            _T_77_44 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_45 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h2d == auto_out_d_bits_source) begin
          _T_77_45 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h2d == auto_in_a_bits_source) begin
              _T_77_45 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h2d == auto_in_a_bits_source) begin
            _T_77_45 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_46 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h2e == auto_out_d_bits_source) begin
          _T_77_46 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h2e == auto_in_a_bits_source) begin
              _T_77_46 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h2e == auto_in_a_bits_source) begin
            _T_77_46 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_47 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h2f == auto_out_d_bits_source) begin
          _T_77_47 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h2f == auto_in_a_bits_source) begin
              _T_77_47 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h2f == auto_in_a_bits_source) begin
            _T_77_47 <= 1'h1;
          end
        end
      end
    end
    if (_T_125) begin
      _T_128 <= _T_32;
    end
    if (reset) begin
      _T_77_48 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h30 == auto_out_d_bits_source) begin
          _T_77_48 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h30 == auto_in_a_bits_source) begin
              _T_77_48 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h30 == auto_in_a_bits_source) begin
            _T_77_48 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_49 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h31 == auto_out_d_bits_source) begin
          _T_77_49 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h31 == auto_in_a_bits_source) begin
              _T_77_49 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h31 == auto_in_a_bits_source) begin
            _T_77_49 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_50 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h32 == auto_out_d_bits_source) begin
          _T_77_50 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h32 == auto_in_a_bits_source) begin
              _T_77_50 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h32 == auto_in_a_bits_source) begin
            _T_77_50 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_51 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h33 == auto_out_d_bits_source) begin
          _T_77_51 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h33 == auto_in_a_bits_source) begin
              _T_77_51 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h33 == auto_in_a_bits_source) begin
            _T_77_51 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_52 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h34 == auto_out_d_bits_source) begin
          _T_77_52 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h34 == auto_in_a_bits_source) begin
              _T_77_52 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h34 == auto_in_a_bits_source) begin
            _T_77_52 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_53 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h35 == auto_out_d_bits_source) begin
          _T_77_53 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h35 == auto_in_a_bits_source) begin
              _T_77_53 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h35 == auto_in_a_bits_source) begin
            _T_77_53 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_54 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h36 == auto_out_d_bits_source) begin
          _T_77_54 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h36 == auto_in_a_bits_source) begin
              _T_77_54 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h36 == auto_in_a_bits_source) begin
            _T_77_54 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_55 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h37 == auto_out_d_bits_source) begin
          _T_77_55 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h37 == auto_in_a_bits_source) begin
              _T_77_55 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h37 == auto_in_a_bits_source) begin
            _T_77_55 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_56 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h38 == auto_out_d_bits_source) begin
          _T_77_56 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h38 == auto_in_a_bits_source) begin
              _T_77_56 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h38 == auto_in_a_bits_source) begin
            _T_77_56 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_57 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h39 == auto_out_d_bits_source) begin
          _T_77_57 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h39 == auto_in_a_bits_source) begin
              _T_77_57 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h39 == auto_in_a_bits_source) begin
            _T_77_57 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_58 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h3a == auto_out_d_bits_source) begin
          _T_77_58 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h3a == auto_in_a_bits_source) begin
              _T_77_58 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h3a == auto_in_a_bits_source) begin
            _T_77_58 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_59 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h3b == auto_out_d_bits_source) begin
          _T_77_59 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h3b == auto_in_a_bits_source) begin
              _T_77_59 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h3b == auto_in_a_bits_source) begin
            _T_77_59 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_60 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h3c == auto_out_d_bits_source) begin
          _T_77_60 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h3c == auto_in_a_bits_source) begin
              _T_77_60 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h3c == auto_in_a_bits_source) begin
            _T_77_60 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_61 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h3d == auto_out_d_bits_source) begin
          _T_77_61 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h3d == auto_in_a_bits_source) begin
              _T_77_61 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h3d == auto_in_a_bits_source) begin
            _T_77_61 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_62 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h3e == auto_out_d_bits_source) begin
          _T_77_62 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h3e == auto_in_a_bits_source) begin
              _T_77_62 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h3e == auto_in_a_bits_source) begin
            _T_77_62 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_63 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h3f == auto_out_d_bits_source) begin
          _T_77_63 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h3f == auto_in_a_bits_source) begin
              _T_77_63 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h3f == auto_in_a_bits_source) begin
            _T_77_63 <= 1'h1;
          end
        end
      end
    end
    if (_T_158) begin
      _T_161 <= _T_32;
    end
    if (reset) begin
      _T_77_64 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h40 == auto_out_d_bits_source) begin
          _T_77_64 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h40 == auto_in_a_bits_source) begin
              _T_77_64 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h40 == auto_in_a_bits_source) begin
            _T_77_64 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_65 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h41 == auto_out_d_bits_source) begin
          _T_77_65 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h41 == auto_in_a_bits_source) begin
              _T_77_65 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h41 == auto_in_a_bits_source) begin
            _T_77_65 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_66 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h42 == auto_out_d_bits_source) begin
          _T_77_66 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h42 == auto_in_a_bits_source) begin
              _T_77_66 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h42 == auto_in_a_bits_source) begin
            _T_77_66 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_67 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h43 == auto_out_d_bits_source) begin
          _T_77_67 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h43 == auto_in_a_bits_source) begin
              _T_77_67 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h43 == auto_in_a_bits_source) begin
            _T_77_67 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_68 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h44 == auto_out_d_bits_source) begin
          _T_77_68 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h44 == auto_in_a_bits_source) begin
              _T_77_68 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h44 == auto_in_a_bits_source) begin
            _T_77_68 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_69 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h45 == auto_out_d_bits_source) begin
          _T_77_69 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h45 == auto_in_a_bits_source) begin
              _T_77_69 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h45 == auto_in_a_bits_source) begin
            _T_77_69 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_70 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h46 == auto_out_d_bits_source) begin
          _T_77_70 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h46 == auto_in_a_bits_source) begin
              _T_77_70 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h46 == auto_in_a_bits_source) begin
            _T_77_70 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_71 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h47 == auto_out_d_bits_source) begin
          _T_77_71 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h47 == auto_in_a_bits_source) begin
              _T_77_71 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h47 == auto_in_a_bits_source) begin
            _T_77_71 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_72 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h48 == auto_out_d_bits_source) begin
          _T_77_72 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h48 == auto_in_a_bits_source) begin
              _T_77_72 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h48 == auto_in_a_bits_source) begin
            _T_77_72 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_73 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h49 == auto_out_d_bits_source) begin
          _T_77_73 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h49 == auto_in_a_bits_source) begin
              _T_77_73 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h49 == auto_in_a_bits_source) begin
            _T_77_73 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_74 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h4a == auto_out_d_bits_source) begin
          _T_77_74 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h4a == auto_in_a_bits_source) begin
              _T_77_74 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h4a == auto_in_a_bits_source) begin
            _T_77_74 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_75 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h4b == auto_out_d_bits_source) begin
          _T_77_75 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h4b == auto_in_a_bits_source) begin
              _T_77_75 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h4b == auto_in_a_bits_source) begin
            _T_77_75 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_76 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h4c == auto_out_d_bits_source) begin
          _T_77_76 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h4c == auto_in_a_bits_source) begin
              _T_77_76 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h4c == auto_in_a_bits_source) begin
            _T_77_76 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_77 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h4d == auto_out_d_bits_source) begin
          _T_77_77 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h4d == auto_in_a_bits_source) begin
              _T_77_77 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h4d == auto_in_a_bits_source) begin
            _T_77_77 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_78 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h4e == auto_out_d_bits_source) begin
          _T_77_78 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h4e == auto_in_a_bits_source) begin
              _T_77_78 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h4e == auto_in_a_bits_source) begin
            _T_77_78 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_79 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h4f == auto_out_d_bits_source) begin
          _T_77_79 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h4f == auto_in_a_bits_source) begin
              _T_77_79 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h4f == auto_in_a_bits_source) begin
            _T_77_79 <= 1'h1;
          end
        end
      end
    end
    if (_T_191) begin
      _T_194 <= _T_32;
    end
    if (reset) begin
      _T_77_80 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h50 == auto_out_d_bits_source) begin
          _T_77_80 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h50 == auto_in_a_bits_source) begin
              _T_77_80 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h50 == auto_in_a_bits_source) begin
            _T_77_80 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_81 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h51 == auto_out_d_bits_source) begin
          _T_77_81 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h51 == auto_in_a_bits_source) begin
              _T_77_81 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h51 == auto_in_a_bits_source) begin
            _T_77_81 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_82 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h52 == auto_out_d_bits_source) begin
          _T_77_82 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h52 == auto_in_a_bits_source) begin
              _T_77_82 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h52 == auto_in_a_bits_source) begin
            _T_77_82 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_83 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h53 == auto_out_d_bits_source) begin
          _T_77_83 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h53 == auto_in_a_bits_source) begin
              _T_77_83 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h53 == auto_in_a_bits_source) begin
            _T_77_83 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_84 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h54 == auto_out_d_bits_source) begin
          _T_77_84 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h54 == auto_in_a_bits_source) begin
              _T_77_84 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h54 == auto_in_a_bits_source) begin
            _T_77_84 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_85 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h55 == auto_out_d_bits_source) begin
          _T_77_85 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h55 == auto_in_a_bits_source) begin
              _T_77_85 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h55 == auto_in_a_bits_source) begin
            _T_77_85 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_86 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h56 == auto_out_d_bits_source) begin
          _T_77_86 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h56 == auto_in_a_bits_source) begin
              _T_77_86 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h56 == auto_in_a_bits_source) begin
            _T_77_86 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_87 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h57 == auto_out_d_bits_source) begin
          _T_77_87 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h57 == auto_in_a_bits_source) begin
              _T_77_87 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h57 == auto_in_a_bits_source) begin
            _T_77_87 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_88 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h58 == auto_out_d_bits_source) begin
          _T_77_88 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h58 == auto_in_a_bits_source) begin
              _T_77_88 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h58 == auto_in_a_bits_source) begin
            _T_77_88 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_89 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h59 == auto_out_d_bits_source) begin
          _T_77_89 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h59 == auto_in_a_bits_source) begin
              _T_77_89 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h59 == auto_in_a_bits_source) begin
            _T_77_89 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_90 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h5a == auto_out_d_bits_source) begin
          _T_77_90 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h5a == auto_in_a_bits_source) begin
              _T_77_90 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h5a == auto_in_a_bits_source) begin
            _T_77_90 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_91 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h5b == auto_out_d_bits_source) begin
          _T_77_91 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h5b == auto_in_a_bits_source) begin
              _T_77_91 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h5b == auto_in_a_bits_source) begin
            _T_77_91 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_92 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h5c == auto_out_d_bits_source) begin
          _T_77_92 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h5c == auto_in_a_bits_source) begin
              _T_77_92 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h5c == auto_in_a_bits_source) begin
            _T_77_92 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_93 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h5d == auto_out_d_bits_source) begin
          _T_77_93 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h5d == auto_in_a_bits_source) begin
              _T_77_93 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h5d == auto_in_a_bits_source) begin
            _T_77_93 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_94 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h5e == auto_out_d_bits_source) begin
          _T_77_94 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h5e == auto_in_a_bits_source) begin
              _T_77_94 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h5e == auto_in_a_bits_source) begin
            _T_77_94 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_95 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h5f == auto_out_d_bits_source) begin
          _T_77_95 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h5f == auto_in_a_bits_source) begin
              _T_77_95 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h5f == auto_in_a_bits_source) begin
            _T_77_95 <= 1'h1;
          end
        end
      end
    end
    if (_T_224) begin
      _T_227 <= _T_32;
    end
    if (reset) begin
      _T_77_96 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h60 == auto_out_d_bits_source) begin
          _T_77_96 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h60 == auto_in_a_bits_source) begin
              _T_77_96 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h60 == auto_in_a_bits_source) begin
            _T_77_96 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_97 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h61 == auto_out_d_bits_source) begin
          _T_77_97 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h61 == auto_in_a_bits_source) begin
              _T_77_97 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h61 == auto_in_a_bits_source) begin
            _T_77_97 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_98 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h62 == auto_out_d_bits_source) begin
          _T_77_98 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h62 == auto_in_a_bits_source) begin
              _T_77_98 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h62 == auto_in_a_bits_source) begin
            _T_77_98 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_99 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h63 == auto_out_d_bits_source) begin
          _T_77_99 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h63 == auto_in_a_bits_source) begin
              _T_77_99 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h63 == auto_in_a_bits_source) begin
            _T_77_99 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_100 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h64 == auto_out_d_bits_source) begin
          _T_77_100 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h64 == auto_in_a_bits_source) begin
              _T_77_100 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h64 == auto_in_a_bits_source) begin
            _T_77_100 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_101 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h65 == auto_out_d_bits_source) begin
          _T_77_101 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h65 == auto_in_a_bits_source) begin
              _T_77_101 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h65 == auto_in_a_bits_source) begin
            _T_77_101 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_102 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h66 == auto_out_d_bits_source) begin
          _T_77_102 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h66 == auto_in_a_bits_source) begin
              _T_77_102 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h66 == auto_in_a_bits_source) begin
            _T_77_102 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_103 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h67 == auto_out_d_bits_source) begin
          _T_77_103 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h67 == auto_in_a_bits_source) begin
              _T_77_103 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h67 == auto_in_a_bits_source) begin
            _T_77_103 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_104 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h68 == auto_out_d_bits_source) begin
          _T_77_104 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h68 == auto_in_a_bits_source) begin
              _T_77_104 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h68 == auto_in_a_bits_source) begin
            _T_77_104 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_105 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h69 == auto_out_d_bits_source) begin
          _T_77_105 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h69 == auto_in_a_bits_source) begin
              _T_77_105 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h69 == auto_in_a_bits_source) begin
            _T_77_105 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_106 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h6a == auto_out_d_bits_source) begin
          _T_77_106 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h6a == auto_in_a_bits_source) begin
              _T_77_106 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h6a == auto_in_a_bits_source) begin
            _T_77_106 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_107 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h6b == auto_out_d_bits_source) begin
          _T_77_107 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h6b == auto_in_a_bits_source) begin
              _T_77_107 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h6b == auto_in_a_bits_source) begin
            _T_77_107 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_108 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h6c == auto_out_d_bits_source) begin
          _T_77_108 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h6c == auto_in_a_bits_source) begin
              _T_77_108 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h6c == auto_in_a_bits_source) begin
            _T_77_108 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_109 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h6d == auto_out_d_bits_source) begin
          _T_77_109 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h6d == auto_in_a_bits_source) begin
              _T_77_109 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h6d == auto_in_a_bits_source) begin
            _T_77_109 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_110 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h6e == auto_out_d_bits_source) begin
          _T_77_110 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h6e == auto_in_a_bits_source) begin
              _T_77_110 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h6e == auto_in_a_bits_source) begin
            _T_77_110 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_111 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h6f == auto_out_d_bits_source) begin
          _T_77_111 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h6f == auto_in_a_bits_source) begin
              _T_77_111 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h6f == auto_in_a_bits_source) begin
            _T_77_111 <= 1'h1;
          end
        end
      end
    end
    if (_T_257) begin
      _T_260 <= _T_32;
    end
    if (reset) begin
      _T_77_112 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h70 == auto_out_d_bits_source) begin
          _T_77_112 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h70 == auto_in_a_bits_source) begin
              _T_77_112 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h70 == auto_in_a_bits_source) begin
            _T_77_112 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_113 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h71 == auto_out_d_bits_source) begin
          _T_77_113 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h71 == auto_in_a_bits_source) begin
              _T_77_113 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h71 == auto_in_a_bits_source) begin
            _T_77_113 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_114 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h72 == auto_out_d_bits_source) begin
          _T_77_114 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h72 == auto_in_a_bits_source) begin
              _T_77_114 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h72 == auto_in_a_bits_source) begin
            _T_77_114 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_115 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h73 == auto_out_d_bits_source) begin
          _T_77_115 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h73 == auto_in_a_bits_source) begin
              _T_77_115 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h73 == auto_in_a_bits_source) begin
            _T_77_115 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_116 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h74 == auto_out_d_bits_source) begin
          _T_77_116 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h74 == auto_in_a_bits_source) begin
              _T_77_116 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h74 == auto_in_a_bits_source) begin
            _T_77_116 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_117 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h75 == auto_out_d_bits_source) begin
          _T_77_117 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h75 == auto_in_a_bits_source) begin
              _T_77_117 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h75 == auto_in_a_bits_source) begin
            _T_77_117 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_118 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h76 == auto_out_d_bits_source) begin
          _T_77_118 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h76 == auto_in_a_bits_source) begin
              _T_77_118 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h76 == auto_in_a_bits_source) begin
            _T_77_118 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_119 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h77 == auto_out_d_bits_source) begin
          _T_77_119 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h77 == auto_in_a_bits_source) begin
              _T_77_119 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h77 == auto_in_a_bits_source) begin
            _T_77_119 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_120 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h78 == auto_out_d_bits_source) begin
          _T_77_120 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h78 == auto_in_a_bits_source) begin
              _T_77_120 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h78 == auto_in_a_bits_source) begin
            _T_77_120 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_121 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h79 == auto_out_d_bits_source) begin
          _T_77_121 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h79 == auto_in_a_bits_source) begin
              _T_77_121 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h79 == auto_in_a_bits_source) begin
            _T_77_121 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_122 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h7a == auto_out_d_bits_source) begin
          _T_77_122 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h7a == auto_in_a_bits_source) begin
              _T_77_122 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h7a == auto_in_a_bits_source) begin
            _T_77_122 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_123 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h7b == auto_out_d_bits_source) begin
          _T_77_123 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h7b == auto_in_a_bits_source) begin
              _T_77_123 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h7b == auto_in_a_bits_source) begin
            _T_77_123 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_124 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h7c == auto_out_d_bits_source) begin
          _T_77_124 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h7c == auto_in_a_bits_source) begin
              _T_77_124 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h7c == auto_in_a_bits_source) begin
            _T_77_124 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_125 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h7d == auto_out_d_bits_source) begin
          _T_77_125 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h7d == auto_in_a_bits_source) begin
              _T_77_125 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h7d == auto_in_a_bits_source) begin
            _T_77_125 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_126 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h7e == auto_out_d_bits_source) begin
          _T_77_126 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h7e == auto_in_a_bits_source) begin
              _T_77_126 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h7e == auto_in_a_bits_source) begin
            _T_77_126 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_77_127 <= 1'h0;
    end else begin
      if (_T_82) begin
        if (7'h7f == auto_out_d_bits_source) begin
          _T_77_127 <= 1'h0;
        end else begin
          if (_T_79) begin
            if (7'h7f == auto_in_a_bits_source) begin
              _T_77_127 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_79) begin
          if (7'h7f == auto_in_a_bits_source) begin
            _T_77_127 <= 1'h1;
          end
        end
      end
    end
    if (_T_290) begin
      _T_293 <= _T_32;
    end
    if (reset) begin
      _T_63 <= 5'h0;
    end else begin
      if (_T_55) begin
        if (_T_66) begin
          if (_T_61) begin
            _T_63 <= _T_60;
          end else begin
            _T_63 <= 5'h0;
          end
        end else begin
          _T_63 <= _T_65;
        end
      end
    end
  end
endmodule
module dual_TLFIFOFixer( 
  input         clock, 
  input         reset, 
  output        auto_in_a_ready, 
  input         auto_in_a_valid, 
  input  [2:0]  auto_in_a_bits_opcode, 
  input  [2:0]  auto_in_a_bits_param, 
  input  [2:0]  auto_in_a_bits_size, 
  input  [2:0]  auto_in_a_bits_source, 
  input  [31:0] auto_in_a_bits_address, 
  input  [3:0]  auto_in_a_bits_mask, 
  input  [31:0] auto_in_a_bits_data, 
  input         auto_in_a_bits_corrupt, 
  input         auto_in_d_ready, 
  output        auto_in_d_valid, 
  output [2:0]  auto_in_d_bits_opcode, 
  output [1:0]  auto_in_d_bits_param, 
  output [2:0]  auto_in_d_bits_size, 
  output [2:0]  auto_in_d_bits_source, 
  output [5:0]  auto_in_d_bits_sink, 
  output        auto_in_d_bits_denied, 
  output [31:0] auto_in_d_bits_data, 
  output        auto_in_d_bits_corrupt, 
  input         auto_out_a_ready, 
  output        auto_out_a_valid, 
  output [2:0]  auto_out_a_bits_opcode, 
  output [2:0]  auto_out_a_bits_param, 
  output [2:0]  auto_out_a_bits_size, 
  output [2:0]  auto_out_a_bits_source, 
  output [31:0] auto_out_a_bits_address, 
  output [3:0]  auto_out_a_bits_mask, 
  output [31:0] auto_out_a_bits_data, 
  output        auto_out_a_bits_corrupt, 
  output        auto_out_d_ready, 
  input         auto_out_d_valid, 
  input  [2:0]  auto_out_d_bits_opcode, 
  input  [1:0]  auto_out_d_bits_param, 
  input  [2:0]  auto_out_d_bits_size, 
  input  [2:0]  auto_out_d_bits_source, 
  input  [5:0]  auto_out_d_bits_sink, 
  input         auto_out_d_bits_denied, 
  input  [31:0] auto_out_d_bits_data, 
  input         auto_out_d_bits_corrupt 
);
  wire  TLMonitor_clock; 
  wire  TLMonitor_reset; 
  wire  TLMonitor_io_in_a_ready; 
  wire  TLMonitor_io_in_a_valid; 
  wire [2:0] TLMonitor_io_in_a_bits_opcode; 
  wire [2:0] TLMonitor_io_in_a_bits_param; 
  wire [2:0] TLMonitor_io_in_a_bits_size; 
  wire [2:0] TLMonitor_io_in_a_bits_source; 
  wire [31:0] TLMonitor_io_in_a_bits_address; 
  wire [3:0] TLMonitor_io_in_a_bits_mask; 
  wire  TLMonitor_io_in_a_bits_corrupt; 
  wire  TLMonitor_io_in_d_ready; 
  wire  TLMonitor_io_in_d_valid; 
  wire [2:0] TLMonitor_io_in_d_bits_opcode; 
  wire [1:0] TLMonitor_io_in_d_bits_param; 
  wire [2:0] TLMonitor_io_in_d_bits_size; 
  wire [2:0] TLMonitor_io_in_d_bits_source; 
  wire [5:0] TLMonitor_io_in_d_bits_sink; 
  wire  TLMonitor_io_in_d_bits_denied; 
  wire  TLMonitor_io_in_d_bits_corrupt; 
  wire [32:0] _T_9; 
  wire [31:0] _T_13; 
  wire [32:0] _T_14; 
  wire [32:0] _T_15; 
  wire [32:0] _T_16; 
  wire  _T_17; 
  wire [31:0] _T_18; 
  wire [32:0] _T_19; 
  wire [32:0] _T_20; 
  wire [32:0] _T_21; 
  wire  _T_22; 
  wire  _T_23; 
  wire [32:0] _T_26; 
  wire [32:0] _T_27; 
  wire  _T_28; 
  wire [1:0] _T_30; 
  wire [1:0] _GEN_38; 
  wire [1:0] _T_31; 
  wire  _T_33; 
  wire  _T_84; 
  wire  _T_85; 
  reg [3:0] _T_43; 
  reg [31:0] _RAND_0;
  wire  _T_46; 
  wire  _T_95; 
  reg  _T_76_0; 
  reg [31:0] _RAND_1;
  reg  _T_76_1; 
  reg [31:0] _RAND_2;
  wire  _T_96; 
  reg  _T_76_2; 
  reg [31:0] _RAND_3;
  wire  _T_97; 
  reg  _T_76_3; 
  reg [31:0] _RAND_4;
  wire  _T_98; 
  wire  _T_99; 
  reg [1:0] _T_94; 
  reg [31:0] _RAND_5;
  wire  _T_100; 
  wire  _T_101; 
  wire  _T_102; 
  wire  _T_116; 
  reg  _T_76_4; 
  reg [31:0] _RAND_6;
  reg  _T_76_5; 
  reg [31:0] _RAND_7;
  wire  _T_117; 
  reg  _T_76_6; 
  reg [31:0] _RAND_8;
  wire  _T_118; 
  reg  _T_76_7; 
  reg [31:0] _RAND_9;
  wire  _T_119; 
  wire  _T_120; 
  reg [1:0] _T_115; 
  reg [31:0] _RAND_10;
  wire  _T_121; 
  wire  _T_122; 
  wire  _T_123; 
  wire  _T_125; 
  wire  _T_129; 
  wire  _T_131; 
  wire  _T_34; 
  wire [12:0] _T_36; 
  wire [5:0] _T_37; 
  wire [5:0] _T_38; 
  wire [3:0] _T_39; 
  wire  _T_40; 
  wire  _T_41; 
  wire [3:0] _T_45; 
  wire  _T_54; 
  wire [12:0] _T_56; 
  wire [5:0] _T_57; 
  wire [5:0] _T_58; 
  wire [3:0] _T_59; 
  wire  _T_60; 
  reg [3:0] _T_62; 
  reg [31:0] _RAND_11;
  wire [3:0] _T_64; 
  wire  _T_65; 
  wire  _T_73; 
  wire  _T_74; 
  wire  _T_78; 
  wire  _T_81; 
  wire  _T_91; 
  wire  _T_112; 
  dual_TLMonitor_11 dual_TLMonitor ( 
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_io_in_a_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt)
  );
  assign _T_9 = {1'b0,$signed(auto_in_a_bits_address)}; 
  assign _T_13 = auto_in_a_bits_address ^ 32'h40000000; 
  assign _T_14 = {1'b0,$signed(_T_13)}; 
  assign _T_15 = $signed(_T_14) & $signed(33'shc0000000); 
  assign _T_16 = $signed(_T_15); 
  assign _T_17 = $signed(_T_16) == $signed(33'sh0); 
  assign _T_18 = auto_in_a_bits_address ^ 32'h80000000; 
  assign _T_19 = {1'b0,$signed(_T_18)}; 
  assign _T_20 = $signed(_T_19) & $signed(33'sh80000000); 
  assign _T_21 = $signed(_T_20); 
  assign _T_22 = $signed(_T_21) == $signed(33'sh0); 
  assign _T_23 = _T_17 | _T_22; 
  assign _T_26 = $signed(_T_9) & $signed(33'shc0000000); 
  assign _T_27 = $signed(_T_26); 
  assign _T_28 = $signed(_T_27) == $signed(33'sh0); 
  assign _T_30 = _T_28 ? 2'h2 : 2'h0; 
  assign _GEN_38 = {{1'd0}, _T_23}; 
  assign _T_31 = _GEN_38 | _T_30; 
  assign _T_33 = _T_31 == 2'h0; 
  assign _T_84 = auto_in_a_bits_source[2:2]; 
  assign _T_85 = _T_84 == 1'h0; 
  assign _T_46 = _T_43 == 4'h0; 
  assign _T_95 = _T_85 & _T_46; 
  assign _T_96 = _T_76_0 | _T_76_1; 
  assign _T_97 = _T_96 | _T_76_2; 
  assign _T_98 = _T_97 | _T_76_3; 
  assign _T_99 = _T_95 & _T_98; 
  assign _T_100 = _T_94 != _T_31; 
  assign _T_101 = _T_33 | _T_100; 
  assign _T_102 = _T_99 & _T_101; 
  assign _T_116 = _T_84 & _T_46; 
  assign _T_117 = _T_76_4 | _T_76_5; 
  assign _T_118 = _T_117 | _T_76_6; 
  assign _T_119 = _T_118 | _T_76_7; 
  assign _T_120 = _T_116 & _T_119; 
  assign _T_121 = _T_115 != _T_31; 
  assign _T_122 = _T_33 | _T_121; 
  assign _T_123 = _T_120 & _T_122; 
  assign _T_125 = _T_102 | _T_123; 
  assign _T_129 = _T_125 == 1'h0; 
  assign _T_131 = auto_out_a_ready & _T_129; 
  assign _T_34 = _T_131 & auto_in_a_valid; 
  assign _T_36 = 13'h3f << auto_in_a_bits_size; 
  assign _T_37 = _T_36[5:0]; 
  assign _T_38 = ~ _T_37; 
  assign _T_39 = _T_38[5:2]; 
  assign _T_40 = auto_in_a_bits_opcode[2]; 
  assign _T_41 = _T_40 == 1'h0; 
  assign _T_45 = _T_43 - 4'h1; 
  assign _T_54 = auto_in_d_ready & auto_out_d_valid; 
  assign _T_56 = 13'h3f << auto_out_d_bits_size; 
  assign _T_57 = _T_56[5:0]; 
  assign _T_58 = ~ _T_57; 
  assign _T_59 = _T_58[5:2]; 
  assign _T_60 = auto_out_d_bits_opcode[0]; 
  assign _T_64 = _T_62 - 4'h1; 
  assign _T_65 = _T_62 == 4'h0; 
  assign _T_73 = auto_out_d_bits_opcode != 3'h6; 
  assign _T_74 = _T_65 & _T_73; 
  assign _T_78 = _T_46 & _T_34; 
  assign _T_81 = _T_74 & _T_54; 
  assign _T_91 = _T_34 & _T_85; 
  assign _T_112 = _T_34 & _T_84; 
  assign auto_in_a_ready = auto_out_a_ready & _T_129; 
  assign auto_in_d_valid = auto_out_d_valid; 
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; 
  assign auto_in_d_bits_param = auto_out_d_bits_param; 
  assign auto_in_d_bits_size = auto_out_d_bits_size; 
  assign auto_in_d_bits_source = auto_out_d_bits_source; 
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; 
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; 
  assign auto_in_d_bits_data = auto_out_d_bits_data; 
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; 
  assign auto_out_a_valid = auto_in_a_valid & _T_129; 
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; 
  assign auto_out_a_bits_param = auto_in_a_bits_param; 
  assign auto_out_a_bits_size = auto_in_a_bits_size; 
  assign auto_out_a_bits_source = auto_in_a_bits_source; 
  assign auto_out_a_bits_address = auto_in_a_bits_address; 
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; 
  assign auto_out_a_bits_data = auto_in_a_bits_data; 
  assign auto_out_a_bits_corrupt = auto_in_a_bits_corrupt; 
  assign auto_out_d_ready = auto_in_d_ready; 
  assign TLMonitor_clock = clock; 
  assign TLMonitor_reset = reset; 
  assign TLMonitor_io_in_a_ready = auto_out_a_ready & _T_129; 
  assign TLMonitor_io_in_a_valid = auto_in_a_valid; 
  assign TLMonitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; 
  assign TLMonitor_io_in_a_bits_param = auto_in_a_bits_param; 
  assign TLMonitor_io_in_a_bits_size = auto_in_a_bits_size; 
  assign TLMonitor_io_in_a_bits_source = auto_in_a_bits_source; 
  assign TLMonitor_io_in_a_bits_address = auto_in_a_bits_address; 
  assign TLMonitor_io_in_a_bits_mask = auto_in_a_bits_mask; 
  assign TLMonitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; 
  assign TLMonitor_io_in_d_ready = auto_in_d_ready; 
  assign TLMonitor_io_in_d_valid = auto_out_d_valid; 
  assign TLMonitor_io_in_d_bits_opcode = auto_out_d_bits_opcode; 
  assign TLMonitor_io_in_d_bits_param = auto_out_d_bits_param; 
  assign TLMonitor_io_in_d_bits_size = auto_out_d_bits_size; 
  assign TLMonitor_io_in_d_bits_source = auto_out_d_bits_source; 
  assign TLMonitor_io_in_d_bits_sink = auto_out_d_bits_sink; 
  assign TLMonitor_io_in_d_bits_denied = auto_out_d_bits_denied; 
  assign TLMonitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_43 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_76_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_76_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_76_2 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_76_3 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_94 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_76_4 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_76_5 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_76_6 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_76_7 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_115 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_62 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_43 <= 4'h0;
    end else begin
      if (_T_34) begin
        if (_T_46) begin
          if (_T_41) begin
            _T_43 <= _T_39;
          end else begin
            _T_43 <= 4'h0;
          end
        end else begin
          _T_43 <= _T_45;
        end
      end
    end
    if (reset) begin
      _T_76_0 <= 1'h0;
    end else begin
      if (_T_81) begin
        if (3'h0 == auto_out_d_bits_source) begin
          _T_76_0 <= 1'h0;
        end else begin
          if (_T_78) begin
            if (3'h0 == auto_in_a_bits_source) begin
              _T_76_0 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_78) begin
          if (3'h0 == auto_in_a_bits_source) begin
            _T_76_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_76_1 <= 1'h0;
    end else begin
      if (_T_81) begin
        if (3'h1 == auto_out_d_bits_source) begin
          _T_76_1 <= 1'h0;
        end else begin
          if (_T_78) begin
            if (3'h1 == auto_in_a_bits_source) begin
              _T_76_1 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_78) begin
          if (3'h1 == auto_in_a_bits_source) begin
            _T_76_1 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_76_2 <= 1'h0;
    end else begin
      if (_T_81) begin
        if (3'h2 == auto_out_d_bits_source) begin
          _T_76_2 <= 1'h0;
        end else begin
          if (_T_78) begin
            if (3'h2 == auto_in_a_bits_source) begin
              _T_76_2 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_78) begin
          if (3'h2 == auto_in_a_bits_source) begin
            _T_76_2 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_76_3 <= 1'h0;
    end else begin
      if (_T_81) begin
        if (3'h3 == auto_out_d_bits_source) begin
          _T_76_3 <= 1'h0;
        end else begin
          if (_T_78) begin
            if (3'h3 == auto_in_a_bits_source) begin
              _T_76_3 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_78) begin
          if (3'h3 == auto_in_a_bits_source) begin
            _T_76_3 <= 1'h1;
          end
        end
      end
    end
    if (_T_91) begin
      _T_94 <= _T_31;
    end
    if (reset) begin
      _T_76_4 <= 1'h0;
    end else begin
      if (_T_81) begin
        if (3'h4 == auto_out_d_bits_source) begin
          _T_76_4 <= 1'h0;
        end else begin
          if (_T_78) begin
            if (3'h4 == auto_in_a_bits_source) begin
              _T_76_4 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_78) begin
          if (3'h4 == auto_in_a_bits_source) begin
            _T_76_4 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_76_5 <= 1'h0;
    end else begin
      if (_T_81) begin
        if (3'h5 == auto_out_d_bits_source) begin
          _T_76_5 <= 1'h0;
        end else begin
          if (_T_78) begin
            if (3'h5 == auto_in_a_bits_source) begin
              _T_76_5 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_78) begin
          if (3'h5 == auto_in_a_bits_source) begin
            _T_76_5 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_76_6 <= 1'h0;
    end else begin
      if (_T_81) begin
        if (3'h6 == auto_out_d_bits_source) begin
          _T_76_6 <= 1'h0;
        end else begin
          if (_T_78) begin
            if (3'h6 == auto_in_a_bits_source) begin
              _T_76_6 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_78) begin
          if (3'h6 == auto_in_a_bits_source) begin
            _T_76_6 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_76_7 <= 1'h0;
    end else begin
      if (_T_81) begin
        if (3'h7 == auto_out_d_bits_source) begin
          _T_76_7 <= 1'h0;
        end else begin
          if (_T_78) begin
            if (3'h7 == auto_in_a_bits_source) begin
              _T_76_7 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_78) begin
          if (3'h7 == auto_in_a_bits_source) begin
            _T_76_7 <= 1'h1;
          end
        end
      end
    end
    if (_T_112) begin
      _T_115 <= _T_31;
    end
    if (reset) begin
      _T_62 <= 4'h0;
    end else begin
      if (_T_54) begin
        if (_T_65) begin
          if (_T_60) begin
            _T_62 <= _T_59;
          end else begin
            _T_62 <= 4'h0;
          end
        end else begin
          _T_62 <= _T_64;
        end
      end
    end
  end
endmodule
module dual_TLHintHandler( 
  input         clock, 
  input         reset, 
  output        auto_in_a_ready, 
  input         auto_in_a_valid, 
  input  [2:0]  auto_in_a_bits_opcode, 
  input  [2:0]  auto_in_a_bits_param, 
  input  [3:0]  auto_in_a_bits_size, 
  input  [5:0]  auto_in_a_bits_source, 
  input  [31:0] auto_in_a_bits_address, 
  input  [7:0]  auto_in_a_bits_mask, 
  input  [63:0] auto_in_a_bits_data, 
  output        auto_in_c_ready, 
  input         auto_in_c_valid, 
  input  [2:0]  auto_in_c_bits_opcode, 
  input  [2:0]  auto_in_c_bits_param, 
  input  [3:0]  auto_in_c_bits_size, 
  input  [5:0]  auto_in_c_bits_source, 
  input  [31:0] auto_in_c_bits_address, 
  input         auto_in_c_bits_corrupt, 
  input         auto_in_d_ready, 
  output        auto_in_d_valid, 
  output [2:0]  auto_in_d_bits_opcode, 
  output [1:0]  auto_in_d_bits_param, 
  output [3:0]  auto_in_d_bits_size, 
  output [5:0]  auto_in_d_bits_source, 
  output        auto_in_d_bits_sink, 
  output        auto_in_d_bits_denied, 
  output [63:0] auto_in_d_bits_data, 
  output        auto_in_d_bits_corrupt, 
  output        auto_in_e_ready, 
  input         auto_in_e_valid, 
  input         auto_in_e_bits_sink, 
  input         auto_out_a_ready, 
  output        auto_out_a_valid, 
  output [2:0]  auto_out_a_bits_opcode, 
  output [2:0]  auto_out_a_bits_param, 
  output [3:0]  auto_out_a_bits_size, 
  output [6:0]  auto_out_a_bits_source, 
  output [31:0] auto_out_a_bits_address, 
  output [7:0]  auto_out_a_bits_mask, 
  output [63:0] auto_out_a_bits_data, 
  input         auto_out_c_ready, 
  output        auto_out_c_valid, 
  output [2:0]  auto_out_c_bits_opcode, 
  output [2:0]  auto_out_c_bits_param, 
  output [3:0]  auto_out_c_bits_size, 
  output [6:0]  auto_out_c_bits_source, 
  output [31:0] auto_out_c_bits_address, 
  output        auto_out_c_bits_corrupt, 
  output        auto_out_d_ready, 
  input         auto_out_d_valid, 
  input  [2:0]  auto_out_d_bits_opcode, 
  input  [1:0]  auto_out_d_bits_param, 
  input  [3:0]  auto_out_d_bits_size, 
  input  [6:0]  auto_out_d_bits_source, 
  input         auto_out_d_bits_sink, 
  input         auto_out_d_bits_denied, 
  input  [63:0] auto_out_d_bits_data, 
  input         auto_out_d_bits_corrupt, 
  input         auto_out_e_ready, 
  output        auto_out_e_valid, 
  output        auto_out_e_bits_sink 
);
  wire  TLMonitor_clock; 
  wire  TLMonitor_reset; 
  wire  TLMonitor_io_in_a_ready; 
  wire  TLMonitor_io_in_a_valid; 
  wire [2:0] TLMonitor_io_in_a_bits_opcode; 
  wire [2:0] TLMonitor_io_in_a_bits_param; 
  wire [3:0] TLMonitor_io_in_a_bits_size; 
  wire [5:0] TLMonitor_io_in_a_bits_source; 
  wire [31:0] TLMonitor_io_in_a_bits_address; 
  wire [7:0] TLMonitor_io_in_a_bits_mask; 
  wire  TLMonitor_io_in_c_ready; 
  wire  TLMonitor_io_in_c_valid; 
  wire [2:0] TLMonitor_io_in_c_bits_opcode; 
  wire [2:0] TLMonitor_io_in_c_bits_param; 
  wire [3:0] TLMonitor_io_in_c_bits_size; 
  wire [5:0] TLMonitor_io_in_c_bits_source; 
  wire [31:0] TLMonitor_io_in_c_bits_address; 
  wire  TLMonitor_io_in_c_bits_corrupt; 
  wire  TLMonitor_io_in_d_ready; 
  wire  TLMonitor_io_in_d_valid; 
  wire [2:0] TLMonitor_io_in_d_bits_opcode; 
  wire [1:0] TLMonitor_io_in_d_bits_param; 
  wire [3:0] TLMonitor_io_in_d_bits_size; 
  wire [5:0] TLMonitor_io_in_d_bits_source; 
  wire  TLMonitor_io_in_d_bits_sink; 
  wire  TLMonitor_io_in_d_bits_denied; 
  wire  TLMonitor_io_in_d_bits_corrupt; 
  wire  TLMonitor_io_in_e_ready; 
  wire  TLMonitor_io_in_e_valid; 
  wire  TLMonitor_io_in_e_bits_sink; 
  wire  Repeater_clock; 
  wire  Repeater_reset; 
  wire  Repeater_io_repeat; 
  wire  Repeater_io_full; 
  wire  Repeater_io_enq_ready; 
  wire  Repeater_io_enq_valid; 
  wire [3:0] Repeater_io_enq_bits_size; 
  wire [5:0] Repeater_io_enq_bits_source; 
  wire [31:0] Repeater_io_enq_bits_address; 
  wire  Repeater_io_deq_ready; 
  wire  Repeater_io_deq_valid; 
  wire [3:0] Repeater_io_deq_bits_size; 
  wire [5:0] Repeater_io_deq_bits_source; 
  wire [31:0] Repeater_io_deq_bits_address; 
  wire  _T_8; 
  wire [31:0] _T_9; 
  wire [32:0] _T_10; 
  wire [32:0] _T_11; 
  wire [32:0] _T_12; 
  wire  _T_13; 
  wire [31:0] _T_14; 
  wire [32:0] _T_15; 
  wire [32:0] _T_16; 
  wire [32:0] _T_17; 
  wire  _T_18; 
  wire  _T_19; 
  wire  _T_29; 
  wire  _T_37_valid; 
  wire  _T_38; 
  wire [3:0] _T_37_bits_size; 
  wire [22:0] _T_40; 
  wire [7:0] _T_41; 
  wire [7:0] _T_42; 
  wire [4:0] _T_43; 
  wire  _T_60; 
  wire [2:0] _T_62; 
  wire  _T_44; 
  wire  _T_45; 
  wire [4:0] _T_46; 
  reg [4:0] _T_47; 
  reg [31:0] _RAND_0;
  wire [4:0] _T_49; 
  wire  _T_50; 
  wire  _T_51; 
  wire  _T_52; 
  wire  _T_53; 
  wire  _T_58; 
  wire [5:0] _T_37_bits_source; 
  wire [6:0] _T_66; 
  wire [6:0] _GEN_1; 
  wire  _T_69; 
  dual_TLMonitor_16 dual_TLMonitor ( 
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_c_ready(TLMonitor_io_in_c_ready),
    .io_in_c_valid(TLMonitor_io_in_c_valid),
    .io_in_c_bits_opcode(TLMonitor_io_in_c_bits_opcode),
    .io_in_c_bits_param(TLMonitor_io_in_c_bits_param),
    .io_in_c_bits_size(TLMonitor_io_in_c_bits_size),
    .io_in_c_bits_source(TLMonitor_io_in_c_bits_source),
    .io_in_c_bits_address(TLMonitor_io_in_c_bits_address),
    .io_in_c_bits_corrupt(TLMonitor_io_in_c_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt),
    .io_in_e_ready(TLMonitor_io_in_e_ready),
    .io_in_e_valid(TLMonitor_io_in_e_valid),
    .io_in_e_bits_sink(TLMonitor_io_in_e_bits_sink)
  );
  dual_Repeater_1 dual_Repeater_top ( 
    .clock(Repeater_clock),
    .reset(Repeater_reset),
    .io_repeat(Repeater_io_repeat),
    .io_full(Repeater_io_full),
    .io_enq_ready(Repeater_io_enq_ready),
    .io_enq_valid(Repeater_io_enq_valid),
    .io_enq_bits_size(Repeater_io_enq_bits_size),
    .io_enq_bits_source(Repeater_io_enq_bits_source),
    .io_enq_bits_address(Repeater_io_enq_bits_address),
    .io_deq_ready(Repeater_io_deq_ready),
    .io_deq_valid(Repeater_io_deq_valid),
    .io_deq_bits_size(Repeater_io_deq_bits_size),
    .io_deq_bits_source(Repeater_io_deq_bits_source),
    .io_deq_bits_address(Repeater_io_deq_bits_address)
  );
  assign _T_8 = auto_in_a_bits_opcode == 3'h5; 
  assign _T_9 = auto_in_a_bits_address ^ 32'h80000000; 
  assign _T_10 = {1'b0,$signed(_T_9)}; 
  assign _T_11 = $signed(_T_10) & $signed(33'sh80000000); 
  assign _T_12 = $signed(_T_11); 
  assign _T_13 = $signed(_T_12) == $signed(33'sh0); 
  assign _T_14 = auto_in_a_bits_address ^ 32'h40000000; 
  assign _T_15 = {1'b0,$signed(_T_14)}; 
  assign _T_16 = $signed(_T_15) & $signed(33'shc0000000); 
  assign _T_17 = $signed(_T_16); 
  assign _T_18 = $signed(_T_17) == $signed(33'sh0); 
  assign _T_19 = _T_13 | _T_18; 
  assign _T_29 = _T_8 & _T_19; 
  assign _T_37_valid = Repeater_io_deq_valid; 
  assign _T_38 = auto_out_a_ready & _T_37_valid; 
  assign _T_37_bits_size = Repeater_io_deq_bits_size; 
  assign _T_40 = 23'hff << _T_37_bits_size; 
  assign _T_41 = _T_40[7:0]; 
  assign _T_42 = ~ _T_41; 
  assign _T_43 = _T_42[7:3]; 
  assign _T_60 = Repeater_io_full | _T_29; 
  assign _T_62 = _T_60 ? 3'h1 : auto_in_a_bits_opcode; 
  assign _T_44 = _T_62[2]; 
  assign _T_45 = _T_44 == 1'h0; 
  assign _T_46 = _T_45 ? _T_43 : 5'h0; 
  assign _T_49 = _T_47 - 5'h1; 
  assign _T_50 = _T_47 == 5'h0; 
  assign _T_51 = _T_47 == 5'h1; 
  assign _T_52 = _T_46 == 5'h0; 
  assign _T_53 = _T_51 | _T_52; 
  assign _T_58 = _T_53 == 1'h0; 
  assign _T_37_bits_source = Repeater_io_deq_bits_source; 
  assign _T_66 = {_T_37_bits_source, 1'h0}; 
  assign _GEN_1 = {{6'd0}, _T_60}; 
  assign _T_69 = auto_out_d_bits_source[0]; 
  assign auto_in_a_ready = Repeater_io_enq_ready; 
  assign auto_in_c_ready = auto_out_c_ready; 
  assign auto_in_d_valid = auto_out_d_valid; 
  assign auto_in_d_bits_opcode = _T_69 ? 3'h2 : auto_out_d_bits_opcode; 
  assign auto_in_d_bits_param = auto_out_d_bits_param; 
  assign auto_in_d_bits_size = auto_out_d_bits_size; 
  assign auto_in_d_bits_source = auto_out_d_bits_source[6:1]; 
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; 
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; 
  assign auto_in_d_bits_data = auto_out_d_bits_data; 
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; 
  assign auto_in_e_ready = auto_out_e_ready; 
  assign auto_out_a_valid = Repeater_io_deq_valid; 
  assign auto_out_a_bits_opcode = _T_60 ? 3'h1 : auto_in_a_bits_opcode; 
  assign auto_out_a_bits_param = _T_60 ? 3'h0 : auto_in_a_bits_param; 
  assign auto_out_a_bits_size = Repeater_io_deq_bits_size; 
  assign auto_out_a_bits_source = _T_66 | _GEN_1; 
  assign auto_out_a_bits_address = Repeater_io_deq_bits_address; 
  assign auto_out_a_bits_mask = _T_60 ? 8'h0 : auto_in_a_bits_mask; 
  assign auto_out_a_bits_data = auto_in_a_bits_data; 
  assign auto_out_c_valid = auto_in_c_valid; 
  assign auto_out_c_bits_opcode = auto_in_c_bits_opcode; 
  assign auto_out_c_bits_param = auto_in_c_bits_param; 
  assign auto_out_c_bits_size = auto_in_c_bits_size; 
  assign auto_out_c_bits_source = {auto_in_c_bits_source, 1'h0}; 
  assign auto_out_c_bits_address = auto_in_c_bits_address; 
  assign auto_out_c_bits_corrupt = auto_in_c_bits_corrupt; 
  assign auto_out_d_ready = auto_in_d_ready; 
  assign auto_out_e_valid = auto_in_e_valid; 
  assign auto_out_e_bits_sink = auto_in_e_bits_sink; 
  assign TLMonitor_clock = clock; 
  assign TLMonitor_reset = reset; 
  assign TLMonitor_io_in_a_ready = Repeater_io_enq_ready; 
  assign TLMonitor_io_in_a_valid = auto_in_a_valid; 
  assign TLMonitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; 
  assign TLMonitor_io_in_a_bits_param = auto_in_a_bits_param; 
  assign TLMonitor_io_in_a_bits_size = auto_in_a_bits_size; 
  assign TLMonitor_io_in_a_bits_source = auto_in_a_bits_source; 
  assign TLMonitor_io_in_a_bits_address = auto_in_a_bits_address; 
  assign TLMonitor_io_in_a_bits_mask = auto_in_a_bits_mask; 
  assign TLMonitor_io_in_c_ready = auto_out_c_ready; 
  assign TLMonitor_io_in_c_valid = auto_in_c_valid; 
  assign TLMonitor_io_in_c_bits_opcode = auto_in_c_bits_opcode; 
  assign TLMonitor_io_in_c_bits_param = auto_in_c_bits_param; 
  assign TLMonitor_io_in_c_bits_size = auto_in_c_bits_size; 
  assign TLMonitor_io_in_c_bits_source = auto_in_c_bits_source; 
  assign TLMonitor_io_in_c_bits_address = auto_in_c_bits_address; 
  assign TLMonitor_io_in_c_bits_corrupt = auto_in_c_bits_corrupt; 
  assign TLMonitor_io_in_d_ready = auto_in_d_ready; 
  assign TLMonitor_io_in_d_valid = auto_out_d_valid; 
  assign TLMonitor_io_in_d_bits_opcode = _T_69 ? 3'h2 : auto_out_d_bits_opcode; 
  assign TLMonitor_io_in_d_bits_param = auto_out_d_bits_param; 
  assign TLMonitor_io_in_d_bits_size = auto_out_d_bits_size; 
  assign TLMonitor_io_in_d_bits_source = auto_out_d_bits_source[6:1]; 
  assign TLMonitor_io_in_d_bits_sink = auto_out_d_bits_sink; 
  assign TLMonitor_io_in_d_bits_denied = auto_out_d_bits_denied; 
  assign TLMonitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; 
  assign TLMonitor_io_in_e_ready = auto_out_e_ready; 
  assign TLMonitor_io_in_e_valid = auto_in_e_valid; 
  assign TLMonitor_io_in_e_bits_sink = auto_in_e_bits_sink; 
  assign Repeater_clock = clock; 
  assign Repeater_reset = reset; 
  assign Repeater_io_repeat = _T_60 & _T_58; 
  assign Repeater_io_enq_valid = auto_in_a_valid; 
  assign Repeater_io_enq_bits_size = auto_in_a_bits_size; 
  assign Repeater_io_enq_bits_source = auto_in_a_bits_source; 
  assign Repeater_io_enq_bits_address = auto_in_a_bits_address; 
  assign Repeater_io_deq_ready = auto_out_a_ready; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_47 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_47 <= 5'h0;
    end else begin
      if (_T_38) begin
        if (_T_50) begin
          if (_T_45) begin
            _T_47 <= _T_43;
          end else begin
            _T_47 <= 5'h0;
          end
        end else begin
          _T_47 <= _T_49;
        end
      end
    end
  end
endmodule
module dual_TLMonitor_10( 
  input         clock, 
  input         reset, 
  input         io_in_a_ready, 
  input         io_in_a_valid, 
  input  [2:0]  io_in_a_bits_opcode, 
  input  [2:0]  io_in_a_bits_param, 
  input  [3:0]  io_in_a_bits_size, 
  input  [6:0]  io_in_a_bits_source, 
  input  [30:0] io_in_a_bits_address, 
  input  [7:0]  io_in_a_bits_mask, 
  input         io_in_a_bits_corrupt, 
  input         io_in_d_ready, 
  input         io_in_d_valid, 
  input  [2:0]  io_in_d_bits_opcode, 
  input  [3:0]  io_in_d_bits_size, 
  input  [6:0]  io_in_d_bits_source, 
  input         io_in_d_bits_denied, 
  input         io_in_d_bits_corrupt 
);
  wire [31:0] plusarg_reader_out; 
  wire [2:0] _T_7; 
  wire  _T_8; 
  wire  _T_16; 
  wire  _T_24; 
  wire  _T_32; 
  wire  _T_40; 
  wire  _T_48; 
  wire  _T_56; 
  wire  _T_64; 
  wire  _T_70; 
  wire  _T_71; 
  wire  _T_72; 
  wire  _T_73; 
  wire  _T_74; 
  wire  _T_75; 
  wire  _T_76; 
  wire [22:0] _T_78; 
  wire [7:0] _T_79; 
  wire [7:0] _T_80; 
  wire [30:0] _GEN_18; 
  wire [30:0] _T_81; 
  wire  _T_82; 
  wire [1:0] _T_84; 
  wire [3:0] _T_85; 
  wire [2:0] _T_86; 
  wire [2:0] _T_87; 
  wire  _T_88; 
  wire  _T_89; 
  wire  _T_90; 
  wire  _T_91; 
  wire  _T_93; 
  wire  _T_94; 
  wire  _T_96; 
  wire  _T_97; 
  wire  _T_98; 
  wire  _T_99; 
  wire  _T_100; 
  wire  _T_101; 
  wire  _T_102; 
  wire  _T_103; 
  wire  _T_104; 
  wire  _T_105; 
  wire  _T_106; 
  wire  _T_107; 
  wire  _T_108; 
  wire  _T_109; 
  wire  _T_110; 
  wire  _T_111; 
  wire  _T_112; 
  wire  _T_113; 
  wire  _T_114; 
  wire  _T_115; 
  wire  _T_116; 
  wire  _T_117; 
  wire  _T_118; 
  wire  _T_119; 
  wire  _T_120; 
  wire  _T_121; 
  wire  _T_122; 
  wire  _T_123; 
  wire  _T_124; 
  wire  _T_125; 
  wire  _T_126; 
  wire  _T_127; 
  wire  _T_128; 
  wire  _T_129; 
  wire  _T_130; 
  wire  _T_131; 
  wire  _T_132; 
  wire  _T_133; 
  wire  _T_134; 
  wire  _T_135; 
  wire  _T_136; 
  wire  _T_137; 
  wire  _T_138; 
  wire  _T_139; 
  wire [7:0] _T_146; 
  wire  _T_277; 
  wire [30:0] _T_279; 
  wire [31:0] _T_280; 
  wire [31:0] _T_281; 
  wire [31:0] _T_282; 
  wire  _T_283; 
  wire  _T_288; 
  wire  _T_355; 
  wire  _T_357; 
  wire  _T_374; 
  wire  _T_375; 
  wire  _T_377; 
  wire  _T_378; 
  wire  _T_381; 
  wire  _T_382; 
  wire  _T_384; 
  wire  _T_385; 
  wire  _T_386; 
  wire  _T_388; 
  wire  _T_389; 
  wire [7:0] _T_390; 
  wire  _T_391; 
  wire  _T_393; 
  wire  _T_394; 
  wire  _T_395; 
  wire  _T_397; 
  wire  _T_398; 
  wire  _T_399; 
  wire  _T_512; 
  wire  _T_514; 
  wire  _T_515; 
  wire  _T_525; 
  wire  _T_535; 
  wire  _T_538; 
  wire  _T_539; 
  wire  _T_546; 
  wire  _T_548; 
  wire  _T_549; 
  wire  _T_550; 
  wire  _T_552; 
  wire  _T_553; 
  wire  _T_558; 
  wire  _T_560; 
  wire  _T_568; 
  wire  _T_571; 
  wire  _T_572; 
  wire  _T_587; 
  wire [7:0] _T_612; 
  wire [7:0] _T_613; 
  wire  _T_614; 
  wire  _T_616; 
  wire  _T_617; 
  wire  _T_618; 
  wire  _T_636; 
  wire  _T_638; 
  wire  _T_639; 
  wire  _T_644; 
  wire  _T_662; 
  wire  _T_664; 
  wire  _T_665; 
  wire  _T_670; 
  wire  _T_696; 
  wire  _T_698; 
  wire  _T_699; 
  wire [2:0] _T_702; 
  wire  _T_703; 
  wire  _T_711; 
  wire  _T_719; 
  wire  _T_727; 
  wire  _T_735; 
  wire  _T_743; 
  wire  _T_751; 
  wire  _T_759; 
  wire  _T_765; 
  wire  _T_766; 
  wire  _T_767; 
  wire  _T_768; 
  wire  _T_769; 
  wire  _T_770; 
  wire  _T_771; 
  wire  _T_773; 
  wire  _T_775; 
  wire  _T_776; 
  wire  _T_777; 
  wire  _T_779; 
  wire  _T_780; 
  wire  _T_785; 
  wire  _T_787; 
  wire  _T_788; 
  wire  _T_789; 
  wire  _T_791; 
  wire  _T_792; 
  wire  _T_793; 
  wire  _T_821; 
  wire  _T_841; 
  wire  _T_843; 
  wire  _T_844; 
  wire  _T_850; 
  wire  _T_867; 
  wire  _T_885; 
  wire  _T_914; 
  wire [4:0] _T_919; 
  wire  _T_920; 
  wire  _T_921; 
  reg [4:0] _T_923; 
  reg [31:0] _RAND_0;
  wire [4:0] _T_925; 
  wire  _T_926; 
  reg [2:0] _T_934; 
  reg [31:0] _RAND_1;
  reg [2:0] _T_935; 
  reg [31:0] _RAND_2;
  reg [3:0] _T_936; 
  reg [31:0] _RAND_3;
  reg [6:0] _T_937; 
  reg [31:0] _RAND_4;
  reg [30:0] _T_938; 
  reg [31:0] _RAND_5;
  wire  _T_939; 
  wire  _T_940; 
  wire  _T_941; 
  wire  _T_943; 
  wire  _T_944; 
  wire  _T_945; 
  wire  _T_947; 
  wire  _T_948; 
  wire  _T_949; 
  wire  _T_951; 
  wire  _T_952; 
  wire  _T_953; 
  wire  _T_955; 
  wire  _T_956; 
  wire  _T_957; 
  wire  _T_959; 
  wire  _T_960; 
  wire  _T_962; 
  wire  _T_963; 
  wire [22:0] _T_965; 
  wire [7:0] _T_966; 
  wire [7:0] _T_967; 
  wire [4:0] _T_968; 
  wire  _T_969; 
  reg [4:0] _T_971; 
  reg [31:0] _RAND_6;
  wire [4:0] _T_973; 
  wire  _T_974; 
  reg [2:0] _T_982; 
  reg [31:0] _RAND_7;
  reg [3:0] _T_984; 
  reg [31:0] _RAND_8;
  reg [6:0] _T_985; 
  reg [31:0] _RAND_9;
  reg  _T_987; 
  reg [31:0] _RAND_10;
  wire  _T_988; 
  wire  _T_989; 
  wire  _T_990; 
  wire  _T_992; 
  wire  _T_993; 
  wire  _T_998; 
  wire  _T_1000; 
  wire  _T_1001; 
  wire  _T_1002; 
  wire  _T_1004; 
  wire  _T_1005; 
  wire  _T_1010; 
  wire  _T_1012; 
  wire  _T_1013; 
  wire  _T_1015; 
  reg [127:0] _T_1016; 
  reg [127:0] _RAND_11;
  reg [4:0] _T_1026; 
  reg [31:0] _RAND_12;
  wire [4:0] _T_1028; 
  wire  _T_1029; 
  reg [4:0] _T_1045; 
  reg [31:0] _RAND_13;
  wire [4:0] _T_1047; 
  wire  _T_1048; 
  wire  _T_1058; 
  wire [127:0] _T_1060; 
  wire [127:0] _T_1061; 
  wire  _T_1062; 
  wire  _T_1063; 
  wire  _T_1065; 
  wire  _T_1066; 
  wire [127:0] _GEN_15; 
  wire  _T_1070; 
  wire  _T_1072; 
  wire  _T_1073; 
  wire [127:0] _T_1074; 
  wire [127:0] _T_1075; 
  wire [127:0] _T_1076; 
  wire  _T_1077; 
  wire  _T_1079; 
  wire  _T_1080; 
  wire [127:0] _GEN_16; 
  wire  _T_1081; 
  wire  _T_1082; 
  wire  _T_1083; 
  wire  _T_1084; 
  wire  _T_1086; 
  wire  _T_1087; 
  wire [127:0] _T_1088; 
  wire [127:0] _T_1089; 
  wire [127:0] _T_1090; 
  reg [31:0] _T_1091; 
  reg [31:0] _RAND_14;
  wire  _T_1092; 
  wire  _T_1093; 
  wire  _T_1094; 
  wire  _T_1095; 
  wire  _T_1096; 
  wire  _T_1097; 
  wire  _T_1099; 
  wire  _T_1100; 
  wire [31:0] _T_1102; 
  wire  _T_1105; 
  wire  _GEN_19; 
  wire  _GEN_35; 
  wire  _GEN_53; 
  wire  _GEN_65; 
  wire  _GEN_75; 
  wire  _GEN_85; 
  wire  _GEN_95; 
  wire  _GEN_105; 
  wire  _GEN_115; 
  wire  _GEN_123; 
  wire  _GEN_131; 
  wire  _GEN_139; 
  wire  _GEN_143; 
  wire  _GEN_147; 
  dual_plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0)) plusarg_reader ( 
    .out(plusarg_reader_out)
  );
  assign _T_7 = io_in_a_bits_source[6:4]; 
  assign _T_8 = _T_7 == 3'h0; 
  assign _T_16 = _T_7 == 3'h1; 
  assign _T_24 = _T_7 == 3'h2; 
  assign _T_32 = _T_7 == 3'h3; 
  assign _T_40 = _T_7 == 3'h4; 
  assign _T_48 = _T_7 == 3'h5; 
  assign _T_56 = _T_7 == 3'h6; 
  assign _T_64 = _T_7 == 3'h7; 
  assign _T_70 = _T_8 | _T_16; 
  assign _T_71 = _T_70 | _T_24; 
  assign _T_72 = _T_71 | _T_32; 
  assign _T_73 = _T_72 | _T_40; 
  assign _T_74 = _T_73 | _T_48; 
  assign _T_75 = _T_74 | _T_56; 
  assign _T_76 = _T_75 | _T_64; 
  assign _T_78 = 23'hff << io_in_a_bits_size; 
  assign _T_79 = _T_78[7:0]; 
  assign _T_80 = ~ _T_79; 
  assign _GEN_18 = {{23'd0}, _T_80}; 
  assign _T_81 = io_in_a_bits_address & _GEN_18; 
  assign _T_82 = _T_81 == 31'h0; 
  assign _T_84 = io_in_a_bits_size[1:0]; 
  assign _T_85 = 4'h1 << _T_84; 
  assign _T_86 = _T_85[2:0]; 
  assign _T_87 = _T_86 | 3'h1; 
  assign _T_88 = io_in_a_bits_size >= 4'h3; 
  assign _T_89 = _T_87[2]; 
  assign _T_90 = io_in_a_bits_address[2]; 
  assign _T_91 = _T_90 == 1'h0; 
  assign _T_93 = _T_89 & _T_91; 
  assign _T_94 = _T_88 | _T_93; 
  assign _T_96 = _T_89 & _T_90; 
  assign _T_97 = _T_88 | _T_96; 
  assign _T_98 = _T_87[1]; 
  assign _T_99 = io_in_a_bits_address[1]; 
  assign _T_100 = _T_99 == 1'h0; 
  assign _T_101 = _T_91 & _T_100; 
  assign _T_102 = _T_98 & _T_101; 
  assign _T_103 = _T_94 | _T_102; 
  assign _T_104 = _T_91 & _T_99; 
  assign _T_105 = _T_98 & _T_104; 
  assign _T_106 = _T_94 | _T_105; 
  assign _T_107 = _T_90 & _T_100; 
  assign _T_108 = _T_98 & _T_107; 
  assign _T_109 = _T_97 | _T_108; 
  assign _T_110 = _T_90 & _T_99; 
  assign _T_111 = _T_98 & _T_110; 
  assign _T_112 = _T_97 | _T_111; 
  assign _T_113 = _T_87[0]; 
  assign _T_114 = io_in_a_bits_address[0]; 
  assign _T_115 = _T_114 == 1'h0; 
  assign _T_116 = _T_101 & _T_115; 
  assign _T_117 = _T_113 & _T_116; 
  assign _T_118 = _T_103 | _T_117; 
  assign _T_119 = _T_101 & _T_114; 
  assign _T_120 = _T_113 & _T_119; 
  assign _T_121 = _T_103 | _T_120; 
  assign _T_122 = _T_104 & _T_115; 
  assign _T_123 = _T_113 & _T_122; 
  assign _T_124 = _T_106 | _T_123; 
  assign _T_125 = _T_104 & _T_114; 
  assign _T_126 = _T_113 & _T_125; 
  assign _T_127 = _T_106 | _T_126; 
  assign _T_128 = _T_107 & _T_115; 
  assign _T_129 = _T_113 & _T_128; 
  assign _T_130 = _T_109 | _T_129; 
  assign _T_131 = _T_107 & _T_114; 
  assign _T_132 = _T_113 & _T_131; 
  assign _T_133 = _T_109 | _T_132; 
  assign _T_134 = _T_110 & _T_115; 
  assign _T_135 = _T_113 & _T_134; 
  assign _T_136 = _T_112 | _T_135; 
  assign _T_137 = _T_110 & _T_114; 
  assign _T_138 = _T_113 & _T_137; 
  assign _T_139 = _T_112 | _T_138; 
  assign _T_146 = {_T_139,_T_136,_T_133,_T_130,_T_127,_T_124,_T_121,_T_118}; 
  assign _T_277 = io_in_a_bits_opcode == 3'h6; 
  assign _T_279 = io_in_a_bits_address ^ 31'h40000000; 
  assign _T_280 = {1'b0,$signed(_T_279)}; 
  assign _T_281 = $signed(_T_280) & $signed(-32'sh20000000); 
  assign _T_282 = $signed(_T_281); 
  assign _T_283 = $signed(_T_282) == $signed(32'sh0); 
  assign _T_288 = reset == 1'h0; 
  assign _T_355 = io_in_a_bits_size <= 4'h6; 
  assign _T_357 = _T_8 ? _T_355 : 1'h0; 
  assign _T_374 = _T_357 | reset; 
  assign _T_375 = _T_374 == 1'h0; 
  assign _T_377 = _T_76 | reset; 
  assign _T_378 = _T_377 == 1'h0; 
  assign _T_381 = _T_88 | reset; 
  assign _T_382 = _T_381 == 1'h0; 
  assign _T_384 = _T_82 | reset; 
  assign _T_385 = _T_384 == 1'h0; 
  assign _T_386 = io_in_a_bits_param <= 3'h2; 
  assign _T_388 = _T_386 | reset; 
  assign _T_389 = _T_388 == 1'h0; 
  assign _T_390 = ~ io_in_a_bits_mask; 
  assign _T_391 = _T_390 == 8'h0; 
  assign _T_393 = _T_391 | reset; 
  assign _T_394 = _T_393 == 1'h0; 
  assign _T_395 = io_in_a_bits_corrupt == 1'h0; 
  assign _T_397 = _T_395 | reset; 
  assign _T_398 = _T_397 == 1'h0; 
  assign _T_399 = io_in_a_bits_opcode == 3'h7; 
  assign _T_512 = io_in_a_bits_param != 3'h0; 
  assign _T_514 = _T_512 | reset; 
  assign _T_515 = _T_514 == 1'h0; 
  assign _T_525 = io_in_a_bits_opcode == 3'h4; 
  assign _T_535 = _T_355 & _T_283; 
  assign _T_538 = _T_535 | reset; 
  assign _T_539 = _T_538 == 1'h0; 
  assign _T_546 = io_in_a_bits_param == 3'h0; 
  assign _T_548 = _T_546 | reset; 
  assign _T_549 = _T_548 == 1'h0; 
  assign _T_550 = io_in_a_bits_mask == _T_146; 
  assign _T_552 = _T_550 | reset; 
  assign _T_553 = _T_552 == 1'h0; 
  assign _T_558 = io_in_a_bits_opcode == 3'h0; 
  assign _T_560 = io_in_a_bits_size <= 4'h8; 
  assign _T_568 = _T_560 & _T_283; 
  assign _T_571 = _T_568 | reset; 
  assign _T_572 = _T_571 == 1'h0; 
  assign _T_587 = io_in_a_bits_opcode == 3'h1; 
  assign _T_612 = ~ _T_146; 
  assign _T_613 = io_in_a_bits_mask & _T_612; 
  assign _T_614 = _T_613 == 8'h0; 
  assign _T_616 = _T_614 | reset; 
  assign _T_617 = _T_616 == 1'h0; 
  assign _T_618 = io_in_a_bits_opcode == 3'h2; 
  assign _T_636 = io_in_a_bits_param <= 3'h4; 
  assign _T_638 = _T_636 | reset; 
  assign _T_639 = _T_638 == 1'h0; 
  assign _T_644 = io_in_a_bits_opcode == 3'h3; 
  assign _T_662 = io_in_a_bits_param <= 3'h3; 
  assign _T_664 = _T_662 | reset; 
  assign _T_665 = _T_664 == 1'h0; 
  assign _T_670 = io_in_a_bits_opcode == 3'h5; 
  assign _T_696 = io_in_d_bits_opcode <= 3'h6; 
  assign _T_698 = _T_696 | reset; 
  assign _T_699 = _T_698 == 1'h0; 
  assign _T_702 = io_in_d_bits_source[6:4]; 
  assign _T_703 = _T_702 == 3'h0; 
  assign _T_711 = _T_702 == 3'h1; 
  assign _T_719 = _T_702 == 3'h2; 
  assign _T_727 = _T_702 == 3'h3; 
  assign _T_735 = _T_702 == 3'h4; 
  assign _T_743 = _T_702 == 3'h5; 
  assign _T_751 = _T_702 == 3'h6; 
  assign _T_759 = _T_702 == 3'h7; 
  assign _T_765 = _T_703 | _T_711; 
  assign _T_766 = _T_765 | _T_719; 
  assign _T_767 = _T_766 | _T_727; 
  assign _T_768 = _T_767 | _T_735; 
  assign _T_769 = _T_768 | _T_743; 
  assign _T_770 = _T_769 | _T_751; 
  assign _T_771 = _T_770 | _T_759; 
  assign _T_773 = io_in_d_bits_opcode == 3'h6; 
  assign _T_775 = _T_771 | reset; 
  assign _T_776 = _T_775 == 1'h0; 
  assign _T_777 = io_in_d_bits_size >= 4'h3; 
  assign _T_779 = _T_777 | reset; 
  assign _T_780 = _T_779 == 1'h0; 
  assign _T_785 = io_in_d_bits_corrupt == 1'h0; 
  assign _T_787 = _T_785 | reset; 
  assign _T_788 = _T_787 == 1'h0; 
  assign _T_789 = io_in_d_bits_denied == 1'h0; 
  assign _T_791 = _T_789 | reset; 
  assign _T_792 = _T_791 == 1'h0; 
  assign _T_793 = io_in_d_bits_opcode == 3'h4; 
  assign _T_821 = io_in_d_bits_opcode == 3'h5; 
  assign _T_841 = _T_789 | io_in_d_bits_corrupt; 
  assign _T_843 = _T_841 | reset; 
  assign _T_844 = _T_843 == 1'h0; 
  assign _T_850 = io_in_d_bits_opcode == 3'h0; 
  assign _T_867 = io_in_d_bits_opcode == 3'h1; 
  assign _T_885 = io_in_d_bits_opcode == 3'h2; 
  assign _T_914 = io_in_a_ready & io_in_a_valid; 
  assign _T_919 = _T_80[7:3]; 
  assign _T_920 = io_in_a_bits_opcode[2]; 
  assign _T_921 = _T_920 == 1'h0; 
  assign _T_925 = _T_923 - 5'h1; 
  assign _T_926 = _T_923 == 5'h0; 
  assign _T_939 = _T_926 == 1'h0; 
  assign _T_940 = io_in_a_valid & _T_939; 
  assign _T_941 = io_in_a_bits_opcode == _T_934; 
  assign _T_943 = _T_941 | reset; 
  assign _T_944 = _T_943 == 1'h0; 
  assign _T_945 = io_in_a_bits_param == _T_935; 
  assign _T_947 = _T_945 | reset; 
  assign _T_948 = _T_947 == 1'h0; 
  assign _T_949 = io_in_a_bits_size == _T_936; 
  assign _T_951 = _T_949 | reset; 
  assign _T_952 = _T_951 == 1'h0; 
  assign _T_953 = io_in_a_bits_source == _T_937; 
  assign _T_955 = _T_953 | reset; 
  assign _T_956 = _T_955 == 1'h0; 
  assign _T_957 = io_in_a_bits_address == _T_938; 
  assign _T_959 = _T_957 | reset; 
  assign _T_960 = _T_959 == 1'h0; 
  assign _T_962 = _T_914 & _T_926; 
  assign _T_963 = io_in_d_ready & io_in_d_valid; 
  assign _T_965 = 23'hff << io_in_d_bits_size; 
  assign _T_966 = _T_965[7:0]; 
  assign _T_967 = ~ _T_966; 
  assign _T_968 = _T_967[7:3]; 
  assign _T_969 = io_in_d_bits_opcode[0]; 
  assign _T_973 = _T_971 - 5'h1; 
  assign _T_974 = _T_971 == 5'h0; 
  assign _T_988 = _T_974 == 1'h0; 
  assign _T_989 = io_in_d_valid & _T_988; 
  assign _T_990 = io_in_d_bits_opcode == _T_982; 
  assign _T_992 = _T_990 | reset; 
  assign _T_993 = _T_992 == 1'h0; 
  assign _T_998 = io_in_d_bits_size == _T_984; 
  assign _T_1000 = _T_998 | reset; 
  assign _T_1001 = _T_1000 == 1'h0; 
  assign _T_1002 = io_in_d_bits_source == _T_985; 
  assign _T_1004 = _T_1002 | reset; 
  assign _T_1005 = _T_1004 == 1'h0; 
  assign _T_1010 = io_in_d_bits_denied == _T_987; 
  assign _T_1012 = _T_1010 | reset; 
  assign _T_1013 = _T_1012 == 1'h0; 
  assign _T_1015 = _T_963 & _T_974; 
  assign _T_1028 = _T_1026 - 5'h1; 
  assign _T_1029 = _T_1026 == 5'h0; 
  assign _T_1047 = _T_1045 - 5'h1; 
  assign _T_1048 = _T_1045 == 5'h0; 
  assign _T_1058 = _T_914 & _T_1029; 
  assign _T_1060 = 128'h1 << io_in_a_bits_source; 
  assign _T_1061 = _T_1016 >> io_in_a_bits_source; 
  assign _T_1062 = _T_1061[0]; 
  assign _T_1063 = _T_1062 == 1'h0; 
  assign _T_1065 = _T_1063 | reset; 
  assign _T_1066 = _T_1065 == 1'h0; 
  assign _GEN_15 = _T_1058 ? _T_1060 : 128'h0; 
  assign _T_1070 = _T_963 & _T_1048; 
  assign _T_1072 = _T_773 == 1'h0; 
  assign _T_1073 = _T_1070 & _T_1072; 
  assign _T_1074 = 128'h1 << io_in_d_bits_source; 
  assign _T_1075 = _GEN_15 | _T_1016; 
  assign _T_1076 = _T_1075 >> io_in_d_bits_source; 
  assign _T_1077 = _T_1076[0]; 
  assign _T_1079 = _T_1077 | reset; 
  assign _T_1080 = _T_1079 == 1'h0; 
  assign _GEN_16 = _T_1073 ? _T_1074 : 128'h0; 
  assign _T_1081 = _GEN_15 != _GEN_16; 
  assign _T_1082 = _GEN_15 != 128'h0; 
  assign _T_1083 = _T_1082 == 1'h0; 
  assign _T_1084 = _T_1081 | _T_1083; 
  assign _T_1086 = _T_1084 | reset; 
  assign _T_1087 = _T_1086 == 1'h0; 
  assign _T_1088 = _T_1016 | _GEN_15; 
  assign _T_1089 = ~ _GEN_16; 
  assign _T_1090 = _T_1088 & _T_1089; 
  assign _T_1092 = _T_1016 != 128'h0; 
  assign _T_1093 = _T_1092 == 1'h0; 
  assign _T_1094 = plusarg_reader_out == 32'h0; 
  assign _T_1095 = _T_1093 | _T_1094; 
  assign _T_1096 = _T_1091 < plusarg_reader_out; 
  assign _T_1097 = _T_1095 | _T_1096; 
  assign _T_1099 = _T_1097 | reset; 
  assign _T_1100 = _T_1099 == 1'h0; 
  assign _T_1102 = _T_1091 + 32'h1; 
  assign _T_1105 = _T_914 | _T_963; 
  assign _GEN_19 = io_in_a_valid & _T_277; 
  assign _GEN_35 = io_in_a_valid & _T_399; 
  assign _GEN_53 = io_in_a_valid & _T_525; 
  assign _GEN_65 = io_in_a_valid & _T_558; 
  assign _GEN_75 = io_in_a_valid & _T_587; 
  assign _GEN_85 = io_in_a_valid & _T_618; 
  assign _GEN_95 = io_in_a_valid & _T_644; 
  assign _GEN_105 = io_in_a_valid & _T_670; 
  assign _GEN_115 = io_in_d_valid & _T_773; 
  assign _GEN_123 = io_in_d_valid & _T_793; 
  assign _GEN_131 = io_in_d_valid & _T_821; 
  assign _GEN_139 = io_in_d_valid & _T_850; 
  assign _GEN_143 = io_in_d_valid & _T_867; 
  assign _GEN_147 = io_in_d_valid & _T_885; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_923 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_934 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_935 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_936 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_937 = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_938 = _RAND_5[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_971 = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_982 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_984 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_985 = _RAND_9[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_987 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {4{`RANDOM}};
  _T_1016 = _RAND_11[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_1026 = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_1045 = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_1091 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_923 <= 5'h0;
    end else begin
      if (_T_914) begin
        if (_T_926) begin
          if (_T_921) begin
            _T_923 <= _T_919;
          end else begin
            _T_923 <= 5'h0;
          end
        end else begin
          _T_923 <= _T_925;
        end
      end
    end
    if (_T_962) begin
      _T_934 <= io_in_a_bits_opcode;
    end
    if (_T_962) begin
      _T_935 <= io_in_a_bits_param;
    end
    if (_T_962) begin
      _T_936 <= io_in_a_bits_size;
    end
    if (_T_962) begin
      _T_937 <= io_in_a_bits_source;
    end
    if (_T_962) begin
      _T_938 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_971 <= 5'h0;
    end else begin
      if (_T_963) begin
        if (_T_974) begin
          if (_T_969) begin
            _T_971 <= _T_968;
          end else begin
            _T_971 <= 5'h0;
          end
        end else begin
          _T_971 <= _T_973;
        end
      end
    end
    if (_T_1015) begin
      _T_982 <= io_in_d_bits_opcode;
    end
    if (_T_1015) begin
      _T_984 <= io_in_d_bits_size;
    end
    if (_T_1015) begin
      _T_985 <= io_in_d_bits_source;
    end
    if (_T_1015) begin
      _T_987 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_1016 <= 128'h0;
    end else begin
      _T_1016 <= _T_1090;
    end
    if (reset) begin
      _T_1026 <= 5'h0;
    end else begin
      if (_T_914) begin
        if (_T_1029) begin
          if (_T_921) begin
            _T_1026 <= _T_919;
          end else begin
            _T_1026 <= 5'h0;
          end
        end else begin
          _T_1026 <= _T_1028;
        end
      end
    end
    if (reset) begin
      _T_1045 <= 5'h0;
    end else begin
      if (_T_963) begin
        if (_T_1048) begin
          if (_T_969) begin
            _T_1045 <= _T_968;
          end else begin
            _T_1045 <= 5'h0;
          end
        end else begin
          _T_1045 <= _T_1047;
        end
      end
    end
    if (reset) begin
      _T_1091 <= 32'h0;
    end else begin
      if (_T_1105) begin
        _T_1091 <= 32'h0;
      end else begin
        _T_1091 <= _T_1102;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel has invalid opcode (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:39 assert (TLMessages.isA(bundle.opcode), \"'A' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:46 assert (visible(edge.address(bundle), bundle.source, edge), \"'A' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_288) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_288) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_375) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_375) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_378) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_378) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_382) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_382) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_385) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_389) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_389) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_394) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_394) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_398) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:56 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_398) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_288) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_288) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_375) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_375) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_378) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_378) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_382) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_382) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_385) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_389) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_389) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_515) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_515) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_394) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_394) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_398) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:68 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_398) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_539) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_539) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_378) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_378) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_385) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_549) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_549) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_553) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_553) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_398) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:77 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_398) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_572) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_572) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_378) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_378) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_385) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_549) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_549) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_553) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_553) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_572) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_572) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_378) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_378) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_385) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_549) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_549) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_617) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_617) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_288) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_288) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_378) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_378) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_385) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_639) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_639) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_553) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_553) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_288) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_288) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_378) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_378) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_385) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_665) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_665) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_553) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_553) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_288) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_288) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_378) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_378) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_385) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_553) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_553) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_398) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:117 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_398) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_699) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_699) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_776) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_776) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_780) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_780) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_788) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_788) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_792) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_792) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_776) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_776) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_288) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:285 assert (sink_ok, \"'D' channel Grant carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_288) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_780) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_780) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_788) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_788) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is denied (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:290 assert (deny_put_ok || !bundle.denied, \"'D' channel Grant is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_776) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_776) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_288) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:295 assert (sink_ok, \"'D' channel GrantData carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_288) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_780) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_780) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_844) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_844) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:300 assert (deny_get_ok || !bundle.denied, \"'D' channel GrantData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_139 & _T_776) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_139 & _T_776) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_139 & _T_788) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_139 & _T_788) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is denied (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:308 assert (deny_put_ok || !bundle.denied, \"'D' channel AccessAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & _T_776) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & _T_776) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & _T_844) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & _T_844) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:316 assert (deny_get_ok || !bundle.denied, \"'D' channel AccessAckData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_147 & _T_776) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_147 & _T_776) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_147 & _T_788) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_147 & _T_788) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is denied (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:324 assert (deny_put_ok || !bundle.denied, \"'D' channel HintAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel valid and not TL-C (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:341 assert (!bundle.b.valid, \"'B' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel valid and not TL-C (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:342 assert (!bundle.c.valid, \"'C' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel valid and not TL-C (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:343 assert (!bundle.e.valid, \"'E' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_940 & _T_944) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_940 & _T_944) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_940 & _T_948) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_940 & _T_948) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_940 & _T_952) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_940 & _T_952) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_940 & _T_956) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_940 & _T_956) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_940 & _T_960) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_940 & _T_960) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_989 & _T_993) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_989 & _T_993) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_989 & _T_1001) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_989 & _T_1001) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_989 & _T_1005) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_989 & _T_1005) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_989 & _T_1013) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_989 & _T_1013) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1058 & _T_1066) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1058 & _T_1066) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1073 & _T_1080) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1073 & _T_1080) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1087) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1087) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1100) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at ChiplinkTest.scala:261:22)\n    at Monitor.scala:479 assert (!inflight.orR || limit === UInt(0) || watchdog < limit, \"TileLink timeout expired\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1100) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLMonitor_11( 
  input         clock, 
  input         reset, 
  input         io_in_a_ready, 
  input         io_in_a_valid, 
  input  [2:0]  io_in_a_bits_opcode, 
  input  [2:0]  io_in_a_bits_param, 
  input  [2:0]  io_in_a_bits_size, 
  input  [2:0]  io_in_a_bits_source, 
  input  [31:0] io_in_a_bits_address, 
  input  [3:0]  io_in_a_bits_mask, 
  input         io_in_a_bits_corrupt, 
  input         io_in_d_ready, 
  input         io_in_d_valid, 
  input  [2:0]  io_in_d_bits_opcode, 
  input  [1:0]  io_in_d_bits_param, 
  input  [2:0]  io_in_d_bits_size, 
  input  [2:0]  io_in_d_bits_source, 
  input  [5:0]  io_in_d_bits_sink, 
  input         io_in_d_bits_denied, 
  input         io_in_d_bits_corrupt 
);
  wire [31:0] plusarg_reader_out; 
  wire  _T_7; 
  wire  _T_8; 
  wire  _T_22; 
  wire [12:0] _T_24; 
  wire [5:0] _T_25; 
  wire [5:0] _T_26; 
  wire [31:0] _GEN_18; 
  wire [31:0] _T_27; 
  wire  _T_28; 
  wire  _T_30; 
  wire [1:0] _T_31; 
  wire [1:0] _T_33; 
  wire  _T_34; 
  wire  _T_35; 
  wire  _T_36; 
  wire  _T_37; 
  wire  _T_39; 
  wire  _T_40; 
  wire  _T_42; 
  wire  _T_43; 
  wire  _T_44; 
  wire  _T_45; 
  wire  _T_46; 
  wire  _T_47; 
  wire  _T_48; 
  wire  _T_49; 
  wire  _T_50; 
  wire  _T_51; 
  wire  _T_52; 
  wire  _T_53; 
  wire  _T_54; 
  wire  _T_55; 
  wire  _T_56; 
  wire  _T_57; 
  wire  _T_58; 
  wire [3:0] _T_61; 
  wire  _T_96; 
  wire [31:0] _T_98; 
  wire [32:0] _T_99; 
  wire [32:0] _T_100; 
  wire [32:0] _T_101; 
  wire  _T_102; 
  wire  _T_104; 
  wire [31:0] _T_106; 
  wire [32:0] _T_107; 
  wire [32:0] _T_108; 
  wire [32:0] _T_109; 
  wire  _T_110; 
  wire  _T_111; 
  wire  _T_113; 
  wire [31:0] _T_116; 
  wire [32:0] _T_117; 
  wire [32:0] _T_118; 
  wire [32:0] _T_119; 
  wire  _T_120; 
  wire  _T_121; 
  wire  _T_124; 
  wire  _T_126; 
  wire  _T_127; 
  wire  _T_130; 
  wire  _T_132; 
  wire  _T_133; 
  wire  _T_136; 
  wire  _T_137; 
  wire  _T_139; 
  wire  _T_140; 
  wire  _T_141; 
  wire  _T_143; 
  wire  _T_144; 
  wire [3:0] _T_145; 
  wire  _T_146; 
  wire  _T_148; 
  wire  _T_149; 
  wire  _T_150; 
  wire  _T_152; 
  wire  _T_153; 
  wire  _T_154; 
  wire  _T_203; 
  wire  _T_205; 
  wire  _T_206; 
  wire  _T_216; 
  wire  _T_236; 
  wire  _T_237; 
  wire  _T_238; 
  wire  _T_241; 
  wire  _T_242; 
  wire  _T_249; 
  wire  _T_251; 
  wire  _T_252; 
  wire  _T_253; 
  wire  _T_255; 
  wire  _T_256; 
  wire  _T_261; 
  wire  _T_302; 
  wire [3:0] _T_339; 
  wire [3:0] _T_340; 
  wire  _T_341; 
  wire  _T_343; 
  wire  _T_344; 
  wire  _T_345; 
  wire  _T_347; 
  wire  _T_361; 
  wire  _T_373; 
  wire  _T_375; 
  wire  _T_376; 
  wire  _T_383; 
  wire  _T_385; 
  wire  _T_386; 
  wire  _T_391; 
  wire  _T_429; 
  wire  _T_431; 
  wire  _T_432; 
  wire  _T_437; 
  wire  _T_478; 
  wire  _T_480; 
  wire  _T_481; 
  wire  _T_484; 
  wire  _T_485; 
  wire  _T_499; 
  wire  _T_500; 
  wire  _T_501; 
  wire  _T_503; 
  wire  _T_504; 
  wire  _T_505; 
  wire  _T_507; 
  wire  _T_508; 
  wire  _T_509; 
  wire  _T_511; 
  wire  _T_512; 
  wire  _T_513; 
  wire  _T_515; 
  wire  _T_516; 
  wire  _T_517; 
  wire  _T_519; 
  wire  _T_520; 
  wire  _T_521; 
  wire  _T_526; 
  wire  _T_527; 
  wire  _T_532; 
  wire  _T_534; 
  wire  _T_535; 
  wire  _T_536; 
  wire  _T_538; 
  wire  _T_539; 
  wire  _T_549; 
  wire  _T_569; 
  wire  _T_571; 
  wire  _T_572; 
  wire  _T_578; 
  wire  _T_595; 
  wire  _T_613; 
  wire  _T_642; 
  wire [3:0] _T_647; 
  wire  _T_648; 
  wire  _T_649; 
  reg [3:0] _T_651; 
  reg [31:0] _RAND_0;
  wire [3:0] _T_653; 
  wire  _T_654; 
  reg [2:0] _T_662; 
  reg [31:0] _RAND_1;
  reg [2:0] _T_663; 
  reg [31:0] _RAND_2;
  reg [2:0] _T_664; 
  reg [31:0] _RAND_3;
  reg [2:0] _T_665; 
  reg [31:0] _RAND_4;
  reg [31:0] _T_666; 
  reg [31:0] _RAND_5;
  wire  _T_667; 
  wire  _T_668; 
  wire  _T_669; 
  wire  _T_671; 
  wire  _T_672; 
  wire  _T_673; 
  wire  _T_675; 
  wire  _T_676; 
  wire  _T_677; 
  wire  _T_679; 
  wire  _T_680; 
  wire  _T_681; 
  wire  _T_683; 
  wire  _T_684; 
  wire  _T_685; 
  wire  _T_687; 
  wire  _T_688; 
  wire  _T_690; 
  wire  _T_691; 
  wire [12:0] _T_693; 
  wire [5:0] _T_694; 
  wire [5:0] _T_695; 
  wire [3:0] _T_696; 
  wire  _T_697; 
  reg [3:0] _T_699; 
  reg [31:0] _RAND_6;
  wire [3:0] _T_701; 
  wire  _T_702; 
  reg [2:0] _T_710; 
  reg [31:0] _RAND_7;
  reg [1:0] _T_711; 
  reg [31:0] _RAND_8;
  reg [2:0] _T_712; 
  reg [31:0] _RAND_9;
  reg [2:0] _T_713; 
  reg [31:0] _RAND_10;
  reg [5:0] _T_714; 
  reg [31:0] _RAND_11;
  reg  _T_715; 
  reg [31:0] _RAND_12;
  wire  _T_716; 
  wire  _T_717; 
  wire  _T_718; 
  wire  _T_720; 
  wire  _T_721; 
  wire  _T_722; 
  wire  _T_724; 
  wire  _T_725; 
  wire  _T_726; 
  wire  _T_728; 
  wire  _T_729; 
  wire  _T_730; 
  wire  _T_732; 
  wire  _T_733; 
  wire  _T_734; 
  wire  _T_736; 
  wire  _T_737; 
  wire  _T_738; 
  wire  _T_740; 
  wire  _T_741; 
  wire  _T_743; 
  reg [7:0] _T_744; 
  reg [31:0] _RAND_13;
  reg [3:0] _T_754; 
  reg [31:0] _RAND_14;
  wire [3:0] _T_756; 
  wire  _T_757; 
  reg [3:0] _T_773; 
  reg [31:0] _RAND_15;
  wire [3:0] _T_775; 
  wire  _T_776; 
  wire  _T_786; 
  wire [7:0] _T_788; 
  wire [7:0] _T_789; 
  wire  _T_790; 
  wire  _T_791; 
  wire  _T_793; 
  wire  _T_794; 
  wire [7:0] _GEN_15; 
  wire  _T_798; 
  wire  _T_800; 
  wire  _T_801; 
  wire [7:0] _T_802; 
  wire [7:0] _T_803; 
  wire [7:0] _T_804; 
  wire  _T_805; 
  wire  _T_807; 
  wire  _T_808; 
  wire [7:0] _GEN_16; 
  wire  _T_809; 
  wire  _T_810; 
  wire  _T_811; 
  wire  _T_812; 
  wire  _T_814; 
  wire  _T_815; 
  wire [7:0] _T_816; 
  wire [7:0] _T_817; 
  wire [7:0] _T_818; 
  reg [31:0] _T_819; 
  reg [31:0] _RAND_16;
  wire  _T_820; 
  wire  _T_821; 
  wire  _T_822; 
  wire  _T_823; 
  wire  _T_824; 
  wire  _T_825; 
  wire  _T_827; 
  wire  _T_828; 
  wire [31:0] _T_830; 
  wire  _T_833; 
  wire  _GEN_19; 
  wire  _GEN_35; 
  wire  _GEN_53; 
  wire  _GEN_65; 
  wire  _GEN_75; 
  wire  _GEN_85; 
  wire  _GEN_95; 
  wire  _GEN_105; 
  wire  _GEN_115; 
  wire  _GEN_125; 
  wire  _GEN_137; 
  wire  _GEN_149; 
  wire  _GEN_155; 
  wire  _GEN_161; 
  dual_plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0)) plusarg_reader ( 
    .out(plusarg_reader_out)
  );
  assign _T_7 = io_in_a_bits_source[2:2]; 
  assign _T_8 = _T_7 == 1'h0; 
  assign _T_22 = _T_8 | _T_7; 
  assign _T_24 = 13'h3f << io_in_a_bits_size; 
  assign _T_25 = _T_24[5:0]; 
  assign _T_26 = ~ _T_25; 
  assign _GEN_18 = {{26'd0}, _T_26}; 
  assign _T_27 = io_in_a_bits_address & _GEN_18; 
  assign _T_28 = _T_27 == 32'h0; 
  assign _T_30 = io_in_a_bits_size[0]; 
  assign _T_31 = 2'h1 << _T_30; 
  assign _T_33 = _T_31 | 2'h1; 
  assign _T_34 = io_in_a_bits_size >= 3'h2; 
  assign _T_35 = _T_33[1]; 
  assign _T_36 = io_in_a_bits_address[1]; 
  assign _T_37 = _T_36 == 1'h0; 
  assign _T_39 = _T_35 & _T_37; 
  assign _T_40 = _T_34 | _T_39; 
  assign _T_42 = _T_35 & _T_36; 
  assign _T_43 = _T_34 | _T_42; 
  assign _T_44 = _T_33[0]; 
  assign _T_45 = io_in_a_bits_address[0]; 
  assign _T_46 = _T_45 == 1'h0; 
  assign _T_47 = _T_37 & _T_46; 
  assign _T_48 = _T_44 & _T_47; 
  assign _T_49 = _T_40 | _T_48; 
  assign _T_50 = _T_37 & _T_45; 
  assign _T_51 = _T_44 & _T_50; 
  assign _T_52 = _T_40 | _T_51; 
  assign _T_53 = _T_36 & _T_46; 
  assign _T_54 = _T_44 & _T_53; 
  assign _T_55 = _T_43 | _T_54; 
  assign _T_56 = _T_36 & _T_45; 
  assign _T_57 = _T_44 & _T_56; 
  assign _T_58 = _T_43 | _T_57; 
  assign _T_61 = {_T_58,_T_55,_T_52,_T_49}; 
  assign _T_96 = io_in_a_bits_opcode == 3'h6; 
  assign _T_98 = io_in_a_bits_address ^ 32'h40000000; 
  assign _T_99 = {1'b0,$signed(_T_98)}; 
  assign _T_100 = $signed(_T_99) & $signed(-33'sh20000000); 
  assign _T_101 = $signed(_T_100); 
  assign _T_102 = $signed(_T_101) == $signed(33'sh0); 
  assign _T_104 = 3'h6 == io_in_a_bits_size; 
  assign _T_106 = io_in_a_bits_address ^ 32'h80000000; 
  assign _T_107 = {1'b0,$signed(_T_106)}; 
  assign _T_108 = $signed(_T_107) & $signed(-33'sh80000000); 
  assign _T_109 = $signed(_T_108); 
  assign _T_110 = $signed(_T_109) == $signed(33'sh0); 
  assign _T_111 = _T_104 & _T_110; 
  assign _T_113 = io_in_a_bits_size <= 3'h6; 
  assign _T_116 = io_in_a_bits_address ^ 32'h10000000; 
  assign _T_117 = {1'b0,$signed(_T_116)}; 
  assign _T_118 = $signed(_T_117) & $signed(-33'sh10000000); 
  assign _T_119 = $signed(_T_118); 
  assign _T_120 = $signed(_T_119) == $signed(33'sh0); 
  assign _T_121 = _T_113 & _T_120; 
  assign _T_124 = _T_111 | _T_121; 
  assign _T_126 = _T_124 | reset; 
  assign _T_127 = _T_126 == 1'h0; 
  assign _T_130 = reset == 1'h0; 
  assign _T_132 = _T_22 | reset; 
  assign _T_133 = _T_132 == 1'h0; 
  assign _T_136 = _T_34 | reset; 
  assign _T_137 = _T_136 == 1'h0; 
  assign _T_139 = _T_28 | reset; 
  assign _T_140 = _T_139 == 1'h0; 
  assign _T_141 = io_in_a_bits_param <= 3'h2; 
  assign _T_143 = _T_141 | reset; 
  assign _T_144 = _T_143 == 1'h0; 
  assign _T_145 = ~ io_in_a_bits_mask; 
  assign _T_146 = _T_145 == 4'h0; 
  assign _T_148 = _T_146 | reset; 
  assign _T_149 = _T_148 == 1'h0; 
  assign _T_150 = io_in_a_bits_corrupt == 1'h0; 
  assign _T_152 = _T_150 | reset; 
  assign _T_153 = _T_152 == 1'h0; 
  assign _T_154 = io_in_a_bits_opcode == 3'h7; 
  assign _T_203 = io_in_a_bits_param != 3'h0; 
  assign _T_205 = _T_203 | reset; 
  assign _T_206 = _T_205 == 1'h0; 
  assign _T_216 = io_in_a_bits_opcode == 3'h4; 
  assign _T_236 = _T_102 | _T_110; 
  assign _T_237 = _T_236 | _T_120; 
  assign _T_238 = _T_113 & _T_237; 
  assign _T_241 = _T_238 | reset; 
  assign _T_242 = _T_241 == 1'h0; 
  assign _T_249 = io_in_a_bits_param == 3'h0; 
  assign _T_251 = _T_249 | reset; 
  assign _T_252 = _T_251 == 1'h0; 
  assign _T_253 = io_in_a_bits_mask == _T_61; 
  assign _T_255 = _T_253 | reset; 
  assign _T_256 = _T_255 == 1'h0; 
  assign _T_261 = io_in_a_bits_opcode == 3'h0; 
  assign _T_302 = io_in_a_bits_opcode == 3'h1; 
  assign _T_339 = ~ _T_61; 
  assign _T_340 = io_in_a_bits_mask & _T_339; 
  assign _T_341 = _T_340 == 4'h0; 
  assign _T_343 = _T_341 | reset; 
  assign _T_344 = _T_343 == 1'h0; 
  assign _T_345 = io_in_a_bits_opcode == 3'h2; 
  assign _T_347 = io_in_a_bits_size <= 3'h3; 
  assign _T_361 = _T_347 & _T_236; 
  assign _T_373 = _T_361 | _T_121; 
  assign _T_375 = _T_373 | reset; 
  assign _T_376 = _T_375 == 1'h0; 
  assign _T_383 = io_in_a_bits_param <= 3'h4; 
  assign _T_385 = _T_383 | reset; 
  assign _T_386 = _T_385 == 1'h0; 
  assign _T_391 = io_in_a_bits_opcode == 3'h3; 
  assign _T_429 = io_in_a_bits_param <= 3'h3; 
  assign _T_431 = _T_429 | reset; 
  assign _T_432 = _T_431 == 1'h0; 
  assign _T_437 = io_in_a_bits_opcode == 3'h5; 
  assign _T_478 = io_in_d_bits_opcode <= 3'h6; 
  assign _T_480 = _T_478 | reset; 
  assign _T_481 = _T_480 == 1'h0; 
  assign _T_484 = io_in_d_bits_source[2:2]; 
  assign _T_485 = _T_484 == 1'h0; 
  assign _T_499 = _T_485 | _T_484; 
  assign _T_500 = io_in_d_bits_sink < 6'h21; 
  assign _T_501 = io_in_d_bits_opcode == 3'h6; 
  assign _T_503 = _T_499 | reset; 
  assign _T_504 = _T_503 == 1'h0; 
  assign _T_505 = io_in_d_bits_size >= 3'h2; 
  assign _T_507 = _T_505 | reset; 
  assign _T_508 = _T_507 == 1'h0; 
  assign _T_509 = io_in_d_bits_param == 2'h0; 
  assign _T_511 = _T_509 | reset; 
  assign _T_512 = _T_511 == 1'h0; 
  assign _T_513 = io_in_d_bits_corrupt == 1'h0; 
  assign _T_515 = _T_513 | reset; 
  assign _T_516 = _T_515 == 1'h0; 
  assign _T_517 = io_in_d_bits_denied == 1'h0; 
  assign _T_519 = _T_517 | reset; 
  assign _T_520 = _T_519 == 1'h0; 
  assign _T_521 = io_in_d_bits_opcode == 3'h4; 
  assign _T_526 = _T_500 | reset; 
  assign _T_527 = _T_526 == 1'h0; 
  assign _T_532 = io_in_d_bits_param <= 2'h2; 
  assign _T_534 = _T_532 | reset; 
  assign _T_535 = _T_534 == 1'h0; 
  assign _T_536 = io_in_d_bits_param != 2'h2; 
  assign _T_538 = _T_536 | reset; 
  assign _T_539 = _T_538 == 1'h0; 
  assign _T_549 = io_in_d_bits_opcode == 3'h5; 
  assign _T_569 = _T_517 | io_in_d_bits_corrupt; 
  assign _T_571 = _T_569 | reset; 
  assign _T_572 = _T_571 == 1'h0; 
  assign _T_578 = io_in_d_bits_opcode == 3'h0; 
  assign _T_595 = io_in_d_bits_opcode == 3'h1; 
  assign _T_613 = io_in_d_bits_opcode == 3'h2; 
  assign _T_642 = io_in_a_ready & io_in_a_valid; 
  assign _T_647 = _T_26[5:2]; 
  assign _T_648 = io_in_a_bits_opcode[2]; 
  assign _T_649 = _T_648 == 1'h0; 
  assign _T_653 = _T_651 - 4'h1; 
  assign _T_654 = _T_651 == 4'h0; 
  assign _T_667 = _T_654 == 1'h0; 
  assign _T_668 = io_in_a_valid & _T_667; 
  assign _T_669 = io_in_a_bits_opcode == _T_662; 
  assign _T_671 = _T_669 | reset; 
  assign _T_672 = _T_671 == 1'h0; 
  assign _T_673 = io_in_a_bits_param == _T_663; 
  assign _T_675 = _T_673 | reset; 
  assign _T_676 = _T_675 == 1'h0; 
  assign _T_677 = io_in_a_bits_size == _T_664; 
  assign _T_679 = _T_677 | reset; 
  assign _T_680 = _T_679 == 1'h0; 
  assign _T_681 = io_in_a_bits_source == _T_665; 
  assign _T_683 = _T_681 | reset; 
  assign _T_684 = _T_683 == 1'h0; 
  assign _T_685 = io_in_a_bits_address == _T_666; 
  assign _T_687 = _T_685 | reset; 
  assign _T_688 = _T_687 == 1'h0; 
  assign _T_690 = _T_642 & _T_654; 
  assign _T_691 = io_in_d_ready & io_in_d_valid; 
  assign _T_693 = 13'h3f << io_in_d_bits_size; 
  assign _T_694 = _T_693[5:0]; 
  assign _T_695 = ~ _T_694; 
  assign _T_696 = _T_695[5:2]; 
  assign _T_697 = io_in_d_bits_opcode[0]; 
  assign _T_701 = _T_699 - 4'h1; 
  assign _T_702 = _T_699 == 4'h0; 
  assign _T_716 = _T_702 == 1'h0; 
  assign _T_717 = io_in_d_valid & _T_716; 
  assign _T_718 = io_in_d_bits_opcode == _T_710; 
  assign _T_720 = _T_718 | reset; 
  assign _T_721 = _T_720 == 1'h0; 
  assign _T_722 = io_in_d_bits_param == _T_711; 
  assign _T_724 = _T_722 | reset; 
  assign _T_725 = _T_724 == 1'h0; 
  assign _T_726 = io_in_d_bits_size == _T_712; 
  assign _T_728 = _T_726 | reset; 
  assign _T_729 = _T_728 == 1'h0; 
  assign _T_730 = io_in_d_bits_source == _T_713; 
  assign _T_732 = _T_730 | reset; 
  assign _T_733 = _T_732 == 1'h0; 
  assign _T_734 = io_in_d_bits_sink == _T_714; 
  assign _T_736 = _T_734 | reset; 
  assign _T_737 = _T_736 == 1'h0; 
  assign _T_738 = io_in_d_bits_denied == _T_715; 
  assign _T_740 = _T_738 | reset; 
  assign _T_741 = _T_740 == 1'h0; 
  assign _T_743 = _T_691 & _T_702; 
  assign _T_756 = _T_754 - 4'h1; 
  assign _T_757 = _T_754 == 4'h0; 
  assign _T_775 = _T_773 - 4'h1; 
  assign _T_776 = _T_773 == 4'h0; 
  assign _T_786 = _T_642 & _T_757; 
  assign _T_788 = 8'h1 << io_in_a_bits_source; 
  assign _T_789 = _T_744 >> io_in_a_bits_source; 
  assign _T_790 = _T_789[0]; 
  assign _T_791 = _T_790 == 1'h0; 
  assign _T_793 = _T_791 | reset; 
  assign _T_794 = _T_793 == 1'h0; 
  assign _GEN_15 = _T_786 ? _T_788 : 8'h0; 
  assign _T_798 = _T_691 & _T_776; 
  assign _T_800 = _T_501 == 1'h0; 
  assign _T_801 = _T_798 & _T_800; 
  assign _T_802 = 8'h1 << io_in_d_bits_source; 
  assign _T_803 = _GEN_15 | _T_744; 
  assign _T_804 = _T_803 >> io_in_d_bits_source; 
  assign _T_805 = _T_804[0]; 
  assign _T_807 = _T_805 | reset; 
  assign _T_808 = _T_807 == 1'h0; 
  assign _GEN_16 = _T_801 ? _T_802 : 8'h0; 
  assign _T_809 = _GEN_15 != _GEN_16; 
  assign _T_810 = _GEN_15 != 8'h0; 
  assign _T_811 = _T_810 == 1'h0; 
  assign _T_812 = _T_809 | _T_811; 
  assign _T_814 = _T_812 | reset; 
  assign _T_815 = _T_814 == 1'h0; 
  assign _T_816 = _T_744 | _GEN_15; 
  assign _T_817 = ~ _GEN_16; 
  assign _T_818 = _T_816 & _T_817; 
  assign _T_820 = _T_744 != 8'h0; 
  assign _T_821 = _T_820 == 1'h0; 
  assign _T_822 = plusarg_reader_out == 32'h0; 
  assign _T_823 = _T_821 | _T_822; 
  assign _T_824 = _T_819 < plusarg_reader_out; 
  assign _T_825 = _T_823 | _T_824; 
  assign _T_827 = _T_825 | reset; 
  assign _T_828 = _T_827 == 1'h0; 
  assign _T_830 = _T_819 + 32'h1; 
  assign _T_833 = _T_642 | _T_691; 
  assign _GEN_19 = io_in_a_valid & _T_96; 
  assign _GEN_35 = io_in_a_valid & _T_154; 
  assign _GEN_53 = io_in_a_valid & _T_216; 
  assign _GEN_65 = io_in_a_valid & _T_261; 
  assign _GEN_75 = io_in_a_valid & _T_302; 
  assign _GEN_85 = io_in_a_valid & _T_345; 
  assign _GEN_95 = io_in_a_valid & _T_391; 
  assign _GEN_105 = io_in_a_valid & _T_437; 
  assign _GEN_115 = io_in_d_valid & _T_501; 
  assign _GEN_125 = io_in_d_valid & _T_521; 
  assign _GEN_137 = io_in_d_valid & _T_549; 
  assign _GEN_149 = io_in_d_valid & _T_578; 
  assign _GEN_155 = io_in_d_valid & _T_595; 
  assign _GEN_161 = io_in_d_valid & _T_613; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_651 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_662 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_663 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_664 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_665 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_666 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_699 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_710 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_711 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_712 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_713 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_714 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_715 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_744 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_754 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_773 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_819 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_651 <= 4'h0;
    end else begin
      if (_T_642) begin
        if (_T_654) begin
          if (_T_649) begin
            _T_651 <= _T_647;
          end else begin
            _T_651 <= 4'h0;
          end
        end else begin
          _T_651 <= _T_653;
        end
      end
    end
    if (_T_690) begin
      _T_662 <= io_in_a_bits_opcode;
    end
    if (_T_690) begin
      _T_663 <= io_in_a_bits_param;
    end
    if (_T_690) begin
      _T_664 <= io_in_a_bits_size;
    end
    if (_T_690) begin
      _T_665 <= io_in_a_bits_source;
    end
    if (_T_690) begin
      _T_666 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_699 <= 4'h0;
    end else begin
      if (_T_691) begin
        if (_T_702) begin
          if (_T_697) begin
            _T_699 <= _T_696;
          end else begin
            _T_699 <= 4'h0;
          end
        end else begin
          _T_699 <= _T_701;
        end
      end
    end
    if (_T_743) begin
      _T_710 <= io_in_d_bits_opcode;
    end
    if (_T_743) begin
      _T_711 <= io_in_d_bits_param;
    end
    if (_T_743) begin
      _T_712 <= io_in_d_bits_size;
    end
    if (_T_743) begin
      _T_713 <= io_in_d_bits_source;
    end
    if (_T_743) begin
      _T_714 <= io_in_d_bits_sink;
    end
    if (_T_743) begin
      _T_715 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_744 <= 8'h0;
    end else begin
      _T_744 <= _T_818;
    end
    if (reset) begin
      _T_754 <= 4'h0;
    end else begin
      if (_T_642) begin
        if (_T_757) begin
          if (_T_649) begin
            _T_754 <= _T_647;
          end else begin
            _T_754 <= 4'h0;
          end
        end else begin
          _T_754 <= _T_756;
        end
      end
    end
    if (reset) begin
      _T_773 <= 4'h0;
    end else begin
      if (_T_691) begin
        if (_T_776) begin
          if (_T_697) begin
            _T_773 <= _T_696;
          end else begin
            _T_773 <= 4'h0;
          end
        end else begin
          _T_773 <= _T_775;
        end
      end
    end
    if (reset) begin
      _T_819 <= 32'h0;
    end else begin
      if (_T_833) begin
        _T_819 <= 32'h0;
      end else begin
        _T_819 <= _T_830;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel has invalid opcode (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:39 assert (TLMessages.isA(bundle.opcode), \"'A' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:46 assert (visible(edge.address(bundle), bundle.source, edge), \"'A' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_127) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_127) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_130) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_130) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_137) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_137) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_140) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_144) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_149) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_149) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_153) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:56 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_153) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_127) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_127) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_130) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_130) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_137) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_137) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_140) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_144) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_206) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_206) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_149) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_149) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_153) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:68 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_153) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_242) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_242) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_140) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_252) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_252) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_256) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_256) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_153) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:77 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_153) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_242) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_242) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_140) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_252) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_252) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_256) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_256) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_242) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_242) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_140) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_252) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_252) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_344) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_344) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_376) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_376) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_140) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_386) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_386) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_256) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_256) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_376) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_376) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_140) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_432) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_432) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_256) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_256) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_242) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_242) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_140) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_256) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_256) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_153) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:117 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_153) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_481) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_481) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_504) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_504) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_508) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_508) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_512) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_512) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_516) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_516) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_520) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_520) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_504) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_504) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_527) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:285 assert (sink_ok, \"'D' channel Grant carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_527) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_508) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_508) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_535) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_535) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_539) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_539) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_516) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_516) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is denied (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:290 assert (deny_put_ok || !bundle.denied, \"'D' channel Grant is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_504) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_504) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_527) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:295 assert (sink_ok, \"'D' channel GrantData carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_527) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_508) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_508) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_535) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_535) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_539) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_539) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_572) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_572) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:300 assert (deny_get_ok || !bundle.denied, \"'D' channel GrantData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_504) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_504) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_512) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_512) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_516) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_516) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is denied (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:308 assert (deny_put_ok || !bundle.denied, \"'D' channel AccessAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_504) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_504) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_512) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_512) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_572) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_572) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:316 assert (deny_get_ok || !bundle.denied, \"'D' channel AccessAckData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_504) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_504) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_512) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_512) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_516) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_516) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is denied (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:324 assert (deny_put_ok || !bundle.denied, \"'D' channel HintAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel valid and not TL-C (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:341 assert (!bundle.b.valid, \"'B' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel valid and not TL-C (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:342 assert (!bundle.c.valid, \"'C' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel valid and not TL-C (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:343 assert (!bundle.e.valid, \"'E' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_668 & _T_672) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_668 & _T_672) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_668 & _T_676) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_668 & _T_676) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_668 & _T_680) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_668 & _T_680) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_668 & _T_684) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_668 & _T_684) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_668 & _T_688) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_668 & _T_688) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_717 & _T_721) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_717 & _T_721) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_717 & _T_725) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_717 & _T_725) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_717 & _T_729) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_717 & _T_729) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_717 & _T_733) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_717 & _T_733) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_717 & _T_737) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_717 & _T_737) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_717 & _T_741) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_717 & _T_741) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_786 & _T_794) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_786 & _T_794) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_801 & _T_808) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_801 & _T_808) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_815) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_815) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_828) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at ChiplinkTest.scala:220:43)\n    at Monitor.scala:479 assert (!inflight.orR || limit === UInt(0) || watchdog < limit, \"TileLink timeout expired\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_828) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLMonitor_12( 
  input         clock, 
  input         reset, 
  input         io_in_a_ready, 
  input         io_in_a_valid, 
  input  [2:0]  io_in_a_bits_opcode, 
  input  [2:0]  io_in_a_bits_param, 
  input  [2:0]  io_in_a_bits_size, 
  input  [2:0]  io_in_a_bits_source, 
  input  [31:0] io_in_a_bits_address, 
  input  [7:0]  io_in_a_bits_mask, 
  input         io_in_a_bits_corrupt, 
  input         io_in_d_ready, 
  input         io_in_d_valid, 
  input  [2:0]  io_in_d_bits_opcode, 
  input  [1:0]  io_in_d_bits_param, 
  input  [2:0]  io_in_d_bits_size, 
  input  [2:0]  io_in_d_bits_source, 
  input  [5:0]  io_in_d_bits_sink, 
  input         io_in_d_bits_denied, 
  input         io_in_d_bits_corrupt 
);
  wire [31:0] plusarg_reader_out; 
  wire  _T_7; 
  wire  _T_8; 
  wire  _T_22; 
  wire [12:0] _T_24; 
  wire [5:0] _T_25; 
  wire [5:0] _T_26; 
  wire [31:0] _GEN_18; 
  wire [31:0] _T_27; 
  wire  _T_28; 
  wire [1:0] _T_30; 
  wire [3:0] _T_31; 
  wire [2:0] _T_32; 
  wire [2:0] _T_33; 
  wire  _T_34; 
  wire  _T_35; 
  wire  _T_36; 
  wire  _T_37; 
  wire  _T_39; 
  wire  _T_40; 
  wire  _T_42; 
  wire  _T_43; 
  wire  _T_44; 
  wire  _T_45; 
  wire  _T_46; 
  wire  _T_47; 
  wire  _T_48; 
  wire  _T_49; 
  wire  _T_50; 
  wire  _T_51; 
  wire  _T_52; 
  wire  _T_53; 
  wire  _T_54; 
  wire  _T_55; 
  wire  _T_56; 
  wire  _T_57; 
  wire  _T_58; 
  wire  _T_59; 
  wire  _T_60; 
  wire  _T_61; 
  wire  _T_62; 
  wire  _T_63; 
  wire  _T_64; 
  wire  _T_65; 
  wire  _T_66; 
  wire  _T_67; 
  wire  _T_68; 
  wire  _T_69; 
  wire  _T_70; 
  wire  _T_71; 
  wire  _T_72; 
  wire  _T_73; 
  wire  _T_74; 
  wire  _T_75; 
  wire  _T_76; 
  wire  _T_77; 
  wire  _T_78; 
  wire  _T_79; 
  wire  _T_80; 
  wire  _T_81; 
  wire  _T_82; 
  wire  _T_83; 
  wire  _T_84; 
  wire  _T_85; 
  wire [7:0] _T_92; 
  wire  _T_127; 
  wire [31:0] _T_129; 
  wire [32:0] _T_130; 
  wire [32:0] _T_131; 
  wire [32:0] _T_132; 
  wire  _T_133; 
  wire  _T_135; 
  wire [31:0] _T_137; 
  wire [32:0] _T_138; 
  wire [32:0] _T_139; 
  wire [32:0] _T_140; 
  wire  _T_141; 
  wire  _T_142; 
  wire  _T_144; 
  wire [31:0] _T_147; 
  wire [32:0] _T_148; 
  wire [32:0] _T_149; 
  wire [32:0] _T_150; 
  wire  _T_151; 
  wire  _T_152; 
  wire  _T_155; 
  wire  _T_157; 
  wire  _T_158; 
  wire  _T_161; 
  wire  _T_163; 
  wire  _T_164; 
  wire  _T_167; 
  wire  _T_168; 
  wire  _T_170; 
  wire  _T_171; 
  wire  _T_172; 
  wire  _T_174; 
  wire  _T_175; 
  wire [7:0] _T_176; 
  wire  _T_177; 
  wire  _T_179; 
  wire  _T_180; 
  wire  _T_181; 
  wire  _T_183; 
  wire  _T_184; 
  wire  _T_185; 
  wire  _T_234; 
  wire  _T_236; 
  wire  _T_237; 
  wire  _T_247; 
  wire  _T_267; 
  wire  _T_268; 
  wire  _T_269; 
  wire  _T_272; 
  wire  _T_273; 
  wire  _T_280; 
  wire  _T_282; 
  wire  _T_283; 
  wire  _T_284; 
  wire  _T_286; 
  wire  _T_287; 
  wire  _T_292; 
  wire  _T_333; 
  wire [7:0] _T_370; 
  wire [7:0] _T_371; 
  wire  _T_372; 
  wire  _T_374; 
  wire  _T_375; 
  wire  _T_376; 
  wire  _T_378; 
  wire  _T_392; 
  wire  _T_404; 
  wire  _T_406; 
  wire  _T_407; 
  wire  _T_414; 
  wire  _T_416; 
  wire  _T_417; 
  wire  _T_422; 
  wire  _T_460; 
  wire  _T_462; 
  wire  _T_463; 
  wire  _T_468; 
  wire  _T_509; 
  wire  _T_511; 
  wire  _T_512; 
  wire  _T_515; 
  wire  _T_516; 
  wire  _T_530; 
  wire  _T_531; 
  wire  _T_532; 
  wire  _T_534; 
  wire  _T_535; 
  wire  _T_536; 
  wire  _T_538; 
  wire  _T_539; 
  wire  _T_540; 
  wire  _T_542; 
  wire  _T_543; 
  wire  _T_544; 
  wire  _T_546; 
  wire  _T_547; 
  wire  _T_548; 
  wire  _T_550; 
  wire  _T_551; 
  wire  _T_552; 
  wire  _T_557; 
  wire  _T_558; 
  wire  _T_563; 
  wire  _T_565; 
  wire  _T_566; 
  wire  _T_567; 
  wire  _T_569; 
  wire  _T_570; 
  wire  _T_580; 
  wire  _T_600; 
  wire  _T_602; 
  wire  _T_603; 
  wire  _T_609; 
  wire  _T_626; 
  wire  _T_644; 
  wire  _T_673; 
  wire [2:0] _T_678; 
  wire  _T_679; 
  wire  _T_680; 
  reg [2:0] _T_682; 
  reg [31:0] _RAND_0;
  wire [2:0] _T_684; 
  wire  _T_685; 
  reg [2:0] _T_693; 
  reg [31:0] _RAND_1;
  reg [2:0] _T_694; 
  reg [31:0] _RAND_2;
  reg [2:0] _T_695; 
  reg [31:0] _RAND_3;
  reg [2:0] _T_696; 
  reg [31:0] _RAND_4;
  reg [31:0] _T_697; 
  reg [31:0] _RAND_5;
  wire  _T_698; 
  wire  _T_699; 
  wire  _T_700; 
  wire  _T_702; 
  wire  _T_703; 
  wire  _T_704; 
  wire  _T_706; 
  wire  _T_707; 
  wire  _T_708; 
  wire  _T_710; 
  wire  _T_711; 
  wire  _T_712; 
  wire  _T_714; 
  wire  _T_715; 
  wire  _T_716; 
  wire  _T_718; 
  wire  _T_719; 
  wire  _T_721; 
  wire  _T_722; 
  wire [12:0] _T_724; 
  wire [5:0] _T_725; 
  wire [5:0] _T_726; 
  wire [2:0] _T_727; 
  wire  _T_728; 
  reg [2:0] _T_730; 
  reg [31:0] _RAND_6;
  wire [2:0] _T_732; 
  wire  _T_733; 
  reg [2:0] _T_741; 
  reg [31:0] _RAND_7;
  reg [1:0] _T_742; 
  reg [31:0] _RAND_8;
  reg [2:0] _T_743; 
  reg [31:0] _RAND_9;
  reg [2:0] _T_744; 
  reg [31:0] _RAND_10;
  reg [5:0] _T_745; 
  reg [31:0] _RAND_11;
  reg  _T_746; 
  reg [31:0] _RAND_12;
  wire  _T_747; 
  wire  _T_748; 
  wire  _T_749; 
  wire  _T_751; 
  wire  _T_752; 
  wire  _T_753; 
  wire  _T_755; 
  wire  _T_756; 
  wire  _T_757; 
  wire  _T_759; 
  wire  _T_760; 
  wire  _T_761; 
  wire  _T_763; 
  wire  _T_764; 
  wire  _T_765; 
  wire  _T_767; 
  wire  _T_768; 
  wire  _T_769; 
  wire  _T_771; 
  wire  _T_772; 
  wire  _T_774; 
  reg [7:0] _T_775; 
  reg [31:0] _RAND_13;
  reg [2:0] _T_785; 
  reg [31:0] _RAND_14;
  wire [2:0] _T_787; 
  wire  _T_788; 
  reg [2:0] _T_804; 
  reg [31:0] _RAND_15;
  wire [2:0] _T_806; 
  wire  _T_807; 
  wire  _T_817; 
  wire [7:0] _T_819; 
  wire [7:0] _T_820; 
  wire  _T_821; 
  wire  _T_822; 
  wire  _T_824; 
  wire  _T_825; 
  wire [7:0] _GEN_15; 
  wire  _T_829; 
  wire  _T_831; 
  wire  _T_832; 
  wire [7:0] _T_833; 
  wire [7:0] _T_834; 
  wire [7:0] _T_835; 
  wire  _T_836; 
  wire  _T_838; 
  wire  _T_839; 
  wire [7:0] _GEN_16; 
  wire  _T_840; 
  wire  _T_841; 
  wire  _T_842; 
  wire  _T_843; 
  wire  _T_845; 
  wire  _T_846; 
  wire [7:0] _T_847; 
  wire [7:0] _T_848; 
  wire [7:0] _T_849; 
  reg [31:0] _T_850; 
  reg [31:0] _RAND_16;
  wire  _T_851; 
  wire  _T_852; 
  wire  _T_853; 
  wire  _T_854; 
  wire  _T_855; 
  wire  _T_856; 
  wire  _T_858; 
  wire  _T_859; 
  wire [31:0] _T_861; 
  wire  _T_864; 
  wire  _GEN_19; 
  wire  _GEN_35; 
  wire  _GEN_53; 
  wire  _GEN_65; 
  wire  _GEN_75; 
  wire  _GEN_85; 
  wire  _GEN_95; 
  wire  _GEN_105; 
  wire  _GEN_115; 
  wire  _GEN_125; 
  wire  _GEN_137; 
  wire  _GEN_149; 
  wire  _GEN_155; 
  wire  _GEN_161; 
  dual_plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0)) plusarg_reader ( 
    .out(plusarg_reader_out)
  );
  assign _T_7 = io_in_a_bits_source[2:2]; 
  assign _T_8 = _T_7 == 1'h0; 
  assign _T_22 = _T_8 | _T_7; 
  assign _T_24 = 13'h3f << io_in_a_bits_size; 
  assign _T_25 = _T_24[5:0]; 
  assign _T_26 = ~ _T_25; 
  assign _GEN_18 = {{26'd0}, _T_26}; 
  assign _T_27 = io_in_a_bits_address & _GEN_18; 
  assign _T_28 = _T_27 == 32'h0; 
  assign _T_30 = io_in_a_bits_size[1:0]; 
  assign _T_31 = 4'h1 << _T_30; 
  assign _T_32 = _T_31[2:0]; 
  assign _T_33 = _T_32 | 3'h1; 
  assign _T_34 = io_in_a_bits_size >= 3'h3; 
  assign _T_35 = _T_33[2]; 
  assign _T_36 = io_in_a_bits_address[2]; 
  assign _T_37 = _T_36 == 1'h0; 
  assign _T_39 = _T_35 & _T_37; 
  assign _T_40 = _T_34 | _T_39; 
  assign _T_42 = _T_35 & _T_36; 
  assign _T_43 = _T_34 | _T_42; 
  assign _T_44 = _T_33[1]; 
  assign _T_45 = io_in_a_bits_address[1]; 
  assign _T_46 = _T_45 == 1'h0; 
  assign _T_47 = _T_37 & _T_46; 
  assign _T_48 = _T_44 & _T_47; 
  assign _T_49 = _T_40 | _T_48; 
  assign _T_50 = _T_37 & _T_45; 
  assign _T_51 = _T_44 & _T_50; 
  assign _T_52 = _T_40 | _T_51; 
  assign _T_53 = _T_36 & _T_46; 
  assign _T_54 = _T_44 & _T_53; 
  assign _T_55 = _T_43 | _T_54; 
  assign _T_56 = _T_36 & _T_45; 
  assign _T_57 = _T_44 & _T_56; 
  assign _T_58 = _T_43 | _T_57; 
  assign _T_59 = _T_33[0]; 
  assign _T_60 = io_in_a_bits_address[0]; 
  assign _T_61 = _T_60 == 1'h0; 
  assign _T_62 = _T_47 & _T_61; 
  assign _T_63 = _T_59 & _T_62; 
  assign _T_64 = _T_49 | _T_63; 
  assign _T_65 = _T_47 & _T_60; 
  assign _T_66 = _T_59 & _T_65; 
  assign _T_67 = _T_49 | _T_66; 
  assign _T_68 = _T_50 & _T_61; 
  assign _T_69 = _T_59 & _T_68; 
  assign _T_70 = _T_52 | _T_69; 
  assign _T_71 = _T_50 & _T_60; 
  assign _T_72 = _T_59 & _T_71; 
  assign _T_73 = _T_52 | _T_72; 
  assign _T_74 = _T_53 & _T_61; 
  assign _T_75 = _T_59 & _T_74; 
  assign _T_76 = _T_55 | _T_75; 
  assign _T_77 = _T_53 & _T_60; 
  assign _T_78 = _T_59 & _T_77; 
  assign _T_79 = _T_55 | _T_78; 
  assign _T_80 = _T_56 & _T_61; 
  assign _T_81 = _T_59 & _T_80; 
  assign _T_82 = _T_58 | _T_81; 
  assign _T_83 = _T_56 & _T_60; 
  assign _T_84 = _T_59 & _T_83; 
  assign _T_85 = _T_58 | _T_84; 
  assign _T_92 = {_T_85,_T_82,_T_79,_T_76,_T_73,_T_70,_T_67,_T_64}; 
  assign _T_127 = io_in_a_bits_opcode == 3'h6; 
  assign _T_129 = io_in_a_bits_address ^ 32'h40000000; 
  assign _T_130 = {1'b0,$signed(_T_129)}; 
  assign _T_131 = $signed(_T_130) & $signed(-33'sh20000000); 
  assign _T_132 = $signed(_T_131); 
  assign _T_133 = $signed(_T_132) == $signed(33'sh0); 
  assign _T_135 = 3'h6 == io_in_a_bits_size; 
  assign _T_137 = io_in_a_bits_address ^ 32'h80000000; 
  assign _T_138 = {1'b0,$signed(_T_137)}; 
  assign _T_139 = $signed(_T_138) & $signed(-33'sh80000000); 
  assign _T_140 = $signed(_T_139); 
  assign _T_141 = $signed(_T_140) == $signed(33'sh0); 
  assign _T_142 = _T_135 & _T_141; 
  assign _T_144 = io_in_a_bits_size <= 3'h6; 
  assign _T_147 = io_in_a_bits_address ^ 32'h10000000; 
  assign _T_148 = {1'b0,$signed(_T_147)}; 
  assign _T_149 = $signed(_T_148) & $signed(-33'sh10000000); 
  assign _T_150 = $signed(_T_149); 
  assign _T_151 = $signed(_T_150) == $signed(33'sh0); 
  assign _T_152 = _T_144 & _T_151; 
  assign _T_155 = _T_142 | _T_152; 
  assign _T_157 = _T_155 | reset; 
  assign _T_158 = _T_157 == 1'h0; 
  assign _T_161 = reset == 1'h0; 
  assign _T_163 = _T_22 | reset; 
  assign _T_164 = _T_163 == 1'h0; 
  assign _T_167 = _T_34 | reset; 
  assign _T_168 = _T_167 == 1'h0; 
  assign _T_170 = _T_28 | reset; 
  assign _T_171 = _T_170 == 1'h0; 
  assign _T_172 = io_in_a_bits_param <= 3'h2; 
  assign _T_174 = _T_172 | reset; 
  assign _T_175 = _T_174 == 1'h0; 
  assign _T_176 = ~ io_in_a_bits_mask; 
  assign _T_177 = _T_176 == 8'h0; 
  assign _T_179 = _T_177 | reset; 
  assign _T_180 = _T_179 == 1'h0; 
  assign _T_181 = io_in_a_bits_corrupt == 1'h0; 
  assign _T_183 = _T_181 | reset; 
  assign _T_184 = _T_183 == 1'h0; 
  assign _T_185 = io_in_a_bits_opcode == 3'h7; 
  assign _T_234 = io_in_a_bits_param != 3'h0; 
  assign _T_236 = _T_234 | reset; 
  assign _T_237 = _T_236 == 1'h0; 
  assign _T_247 = io_in_a_bits_opcode == 3'h4; 
  assign _T_267 = _T_133 | _T_141; 
  assign _T_268 = _T_267 | _T_151; 
  assign _T_269 = _T_144 & _T_268; 
  assign _T_272 = _T_269 | reset; 
  assign _T_273 = _T_272 == 1'h0; 
  assign _T_280 = io_in_a_bits_param == 3'h0; 
  assign _T_282 = _T_280 | reset; 
  assign _T_283 = _T_282 == 1'h0; 
  assign _T_284 = io_in_a_bits_mask == _T_92; 
  assign _T_286 = _T_284 | reset; 
  assign _T_287 = _T_286 == 1'h0; 
  assign _T_292 = io_in_a_bits_opcode == 3'h0; 
  assign _T_333 = io_in_a_bits_opcode == 3'h1; 
  assign _T_370 = ~ _T_92; 
  assign _T_371 = io_in_a_bits_mask & _T_370; 
  assign _T_372 = _T_371 == 8'h0; 
  assign _T_374 = _T_372 | reset; 
  assign _T_375 = _T_374 == 1'h0; 
  assign _T_376 = io_in_a_bits_opcode == 3'h2; 
  assign _T_378 = io_in_a_bits_size <= 3'h3; 
  assign _T_392 = _T_378 & _T_267; 
  assign _T_404 = _T_392 | _T_152; 
  assign _T_406 = _T_404 | reset; 
  assign _T_407 = _T_406 == 1'h0; 
  assign _T_414 = io_in_a_bits_param <= 3'h4; 
  assign _T_416 = _T_414 | reset; 
  assign _T_417 = _T_416 == 1'h0; 
  assign _T_422 = io_in_a_bits_opcode == 3'h3; 
  assign _T_460 = io_in_a_bits_param <= 3'h3; 
  assign _T_462 = _T_460 | reset; 
  assign _T_463 = _T_462 == 1'h0; 
  assign _T_468 = io_in_a_bits_opcode == 3'h5; 
  assign _T_509 = io_in_d_bits_opcode <= 3'h6; 
  assign _T_511 = _T_509 | reset; 
  assign _T_512 = _T_511 == 1'h0; 
  assign _T_515 = io_in_d_bits_source[2:2]; 
  assign _T_516 = _T_515 == 1'h0; 
  assign _T_530 = _T_516 | _T_515; 
  assign _T_531 = io_in_d_bits_sink < 6'h21; 
  assign _T_532 = io_in_d_bits_opcode == 3'h6; 
  assign _T_534 = _T_530 | reset; 
  assign _T_535 = _T_534 == 1'h0; 
  assign _T_536 = io_in_d_bits_size >= 3'h3; 
  assign _T_538 = _T_536 | reset; 
  assign _T_539 = _T_538 == 1'h0; 
  assign _T_540 = io_in_d_bits_param == 2'h0; 
  assign _T_542 = _T_540 | reset; 
  assign _T_543 = _T_542 == 1'h0; 
  assign _T_544 = io_in_d_bits_corrupt == 1'h0; 
  assign _T_546 = _T_544 | reset; 
  assign _T_547 = _T_546 == 1'h0; 
  assign _T_548 = io_in_d_bits_denied == 1'h0; 
  assign _T_550 = _T_548 | reset; 
  assign _T_551 = _T_550 == 1'h0; 
  assign _T_552 = io_in_d_bits_opcode == 3'h4; 
  assign _T_557 = _T_531 | reset; 
  assign _T_558 = _T_557 == 1'h0; 
  assign _T_563 = io_in_d_bits_param <= 2'h2; 
  assign _T_565 = _T_563 | reset; 
  assign _T_566 = _T_565 == 1'h0; 
  assign _T_567 = io_in_d_bits_param != 2'h2; 
  assign _T_569 = _T_567 | reset; 
  assign _T_570 = _T_569 == 1'h0; 
  assign _T_580 = io_in_d_bits_opcode == 3'h5; 
  assign _T_600 = _T_548 | io_in_d_bits_corrupt; 
  assign _T_602 = _T_600 | reset; 
  assign _T_603 = _T_602 == 1'h0; 
  assign _T_609 = io_in_d_bits_opcode == 3'h0; 
  assign _T_626 = io_in_d_bits_opcode == 3'h1; 
  assign _T_644 = io_in_d_bits_opcode == 3'h2; 
  assign _T_673 = io_in_a_ready & io_in_a_valid; 
  assign _T_678 = _T_26[5:3]; 
  assign _T_679 = io_in_a_bits_opcode[2]; 
  assign _T_680 = _T_679 == 1'h0; 
  assign _T_684 = _T_682 - 3'h1; 
  assign _T_685 = _T_682 == 3'h0; 
  assign _T_698 = _T_685 == 1'h0; 
  assign _T_699 = io_in_a_valid & _T_698; 
  assign _T_700 = io_in_a_bits_opcode == _T_693; 
  assign _T_702 = _T_700 | reset; 
  assign _T_703 = _T_702 == 1'h0; 
  assign _T_704 = io_in_a_bits_param == _T_694; 
  assign _T_706 = _T_704 | reset; 
  assign _T_707 = _T_706 == 1'h0; 
  assign _T_708 = io_in_a_bits_size == _T_695; 
  assign _T_710 = _T_708 | reset; 
  assign _T_711 = _T_710 == 1'h0; 
  assign _T_712 = io_in_a_bits_source == _T_696; 
  assign _T_714 = _T_712 | reset; 
  assign _T_715 = _T_714 == 1'h0; 
  assign _T_716 = io_in_a_bits_address == _T_697; 
  assign _T_718 = _T_716 | reset; 
  assign _T_719 = _T_718 == 1'h0; 
  assign _T_721 = _T_673 & _T_685; 
  assign _T_722 = io_in_d_ready & io_in_d_valid; 
  assign _T_724 = 13'h3f << io_in_d_bits_size; 
  assign _T_725 = _T_724[5:0]; 
  assign _T_726 = ~ _T_725; 
  assign _T_727 = _T_726[5:3]; 
  assign _T_728 = io_in_d_bits_opcode[0]; 
  assign _T_732 = _T_730 - 3'h1; 
  assign _T_733 = _T_730 == 3'h0; 
  assign _T_747 = _T_733 == 1'h0; 
  assign _T_748 = io_in_d_valid & _T_747; 
  assign _T_749 = io_in_d_bits_opcode == _T_741; 
  assign _T_751 = _T_749 | reset; 
  assign _T_752 = _T_751 == 1'h0; 
  assign _T_753 = io_in_d_bits_param == _T_742; 
  assign _T_755 = _T_753 | reset; 
  assign _T_756 = _T_755 == 1'h0; 
  assign _T_757 = io_in_d_bits_size == _T_743; 
  assign _T_759 = _T_757 | reset; 
  assign _T_760 = _T_759 == 1'h0; 
  assign _T_761 = io_in_d_bits_source == _T_744; 
  assign _T_763 = _T_761 | reset; 
  assign _T_764 = _T_763 == 1'h0; 
  assign _T_765 = io_in_d_bits_sink == _T_745; 
  assign _T_767 = _T_765 | reset; 
  assign _T_768 = _T_767 == 1'h0; 
  assign _T_769 = io_in_d_bits_denied == _T_746; 
  assign _T_771 = _T_769 | reset; 
  assign _T_772 = _T_771 == 1'h0; 
  assign _T_774 = _T_722 & _T_733; 
  assign _T_787 = _T_785 - 3'h1; 
  assign _T_788 = _T_785 == 3'h0; 
  assign _T_806 = _T_804 - 3'h1; 
  assign _T_807 = _T_804 == 3'h0; 
  assign _T_817 = _T_673 & _T_788; 
  assign _T_819 = 8'h1 << io_in_a_bits_source; 
  assign _T_820 = _T_775 >> io_in_a_bits_source; 
  assign _T_821 = _T_820[0]; 
  assign _T_822 = _T_821 == 1'h0; 
  assign _T_824 = _T_822 | reset; 
  assign _T_825 = _T_824 == 1'h0; 
  assign _GEN_15 = _T_817 ? _T_819 : 8'h0; 
  assign _T_829 = _T_722 & _T_807; 
  assign _T_831 = _T_532 == 1'h0; 
  assign _T_832 = _T_829 & _T_831; 
  assign _T_833 = 8'h1 << io_in_d_bits_source; 
  assign _T_834 = _GEN_15 | _T_775; 
  assign _T_835 = _T_834 >> io_in_d_bits_source; 
  assign _T_836 = _T_835[0]; 
  assign _T_838 = _T_836 | reset; 
  assign _T_839 = _T_838 == 1'h0; 
  assign _GEN_16 = _T_832 ? _T_833 : 8'h0; 
  assign _T_840 = _GEN_15 != _GEN_16; 
  assign _T_841 = _GEN_15 != 8'h0; 
  assign _T_842 = _T_841 == 1'h0; 
  assign _T_843 = _T_840 | _T_842; 
  assign _T_845 = _T_843 | reset; 
  assign _T_846 = _T_845 == 1'h0; 
  assign _T_847 = _T_775 | _GEN_15; 
  assign _T_848 = ~ _GEN_16; 
  assign _T_849 = _T_847 & _T_848; 
  assign _T_851 = _T_775 != 8'h0; 
  assign _T_852 = _T_851 == 1'h0; 
  assign _T_853 = plusarg_reader_out == 32'h0; 
  assign _T_854 = _T_852 | _T_853; 
  assign _T_855 = _T_850 < plusarg_reader_out; 
  assign _T_856 = _T_854 | _T_855; 
  assign _T_858 = _T_856 | reset; 
  assign _T_859 = _T_858 == 1'h0; 
  assign _T_861 = _T_850 + 32'h1; 
  assign _T_864 = _T_673 | _T_722; 
  assign _GEN_19 = io_in_a_valid & _T_127; 
  assign _GEN_35 = io_in_a_valid & _T_185; 
  assign _GEN_53 = io_in_a_valid & _T_247; 
  assign _GEN_65 = io_in_a_valid & _T_292; 
  assign _GEN_75 = io_in_a_valid & _T_333; 
  assign _GEN_85 = io_in_a_valid & _T_376; 
  assign _GEN_95 = io_in_a_valid & _T_422; 
  assign _GEN_105 = io_in_a_valid & _T_468; 
  assign _GEN_115 = io_in_d_valid & _T_532; 
  assign _GEN_125 = io_in_d_valid & _T_552; 
  assign _GEN_137 = io_in_d_valid & _T_580; 
  assign _GEN_149 = io_in_d_valid & _T_609; 
  assign _GEN_155 = io_in_d_valid & _T_626; 
  assign _GEN_161 = io_in_d_valid & _T_644; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_682 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_693 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_694 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_695 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_696 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_697 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_730 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_741 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_742 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_743 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_744 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_745 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_746 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_775 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_785 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_804 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_850 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_682 <= 3'h0;
    end else begin
      if (_T_673) begin
        if (_T_685) begin
          if (_T_680) begin
            _T_682 <= _T_678;
          end else begin
            _T_682 <= 3'h0;
          end
        end else begin
          _T_682 <= _T_684;
        end
      end
    end
    if (_T_721) begin
      _T_693 <= io_in_a_bits_opcode;
    end
    if (_T_721) begin
      _T_694 <= io_in_a_bits_param;
    end
    if (_T_721) begin
      _T_695 <= io_in_a_bits_size;
    end
    if (_T_721) begin
      _T_696 <= io_in_a_bits_source;
    end
    if (_T_721) begin
      _T_697 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_730 <= 3'h0;
    end else begin
      if (_T_722) begin
        if (_T_733) begin
          if (_T_728) begin
            _T_730 <= _T_727;
          end else begin
            _T_730 <= 3'h0;
          end
        end else begin
          _T_730 <= _T_732;
        end
      end
    end
    if (_T_774) begin
      _T_741 <= io_in_d_bits_opcode;
    end
    if (_T_774) begin
      _T_742 <= io_in_d_bits_param;
    end
    if (_T_774) begin
      _T_743 <= io_in_d_bits_size;
    end
    if (_T_774) begin
      _T_744 <= io_in_d_bits_source;
    end
    if (_T_774) begin
      _T_745 <= io_in_d_bits_sink;
    end
    if (_T_774) begin
      _T_746 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_775 <= 8'h0;
    end else begin
      _T_775 <= _T_849;
    end
    if (reset) begin
      _T_785 <= 3'h0;
    end else begin
      if (_T_673) begin
        if (_T_788) begin
          if (_T_680) begin
            _T_785 <= _T_678;
          end else begin
            _T_785 <= 3'h0;
          end
        end else begin
          _T_785 <= _T_787;
        end
      end
    end
    if (reset) begin
      _T_804 <= 3'h0;
    end else begin
      if (_T_722) begin
        if (_T_807) begin
          if (_T_728) begin
            _T_804 <= _T_727;
          end else begin
            _T_804 <= 3'h0;
          end
        end else begin
          _T_804 <= _T_806;
        end
      end
    end
    if (reset) begin
      _T_850 <= 32'h0;
    end else begin
      if (_T_864) begin
        _T_850 <= 32'h0;
      end else begin
        _T_850 <= _T_861;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel has invalid opcode (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:39 assert (TLMessages.isA(bundle.opcode), \"'A' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:46 assert (visible(edge.address(bundle), bundle.source, edge), \"'A' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_158) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_158) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_161) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_161) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_164) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_164) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_168) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_168) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_171) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_171) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_175) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_175) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_180) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_180) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_184) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:56 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_184) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_158) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_158) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_161) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_161) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_164) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_164) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_168) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_168) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_171) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_171) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_175) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_175) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_237) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_237) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_180) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_180) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_184) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:68 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_184) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_273) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_273) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_164) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_164) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_171) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_171) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_283) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_283) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_287) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_287) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_184) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:77 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_184) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_273) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_273) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_164) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_164) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_171) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_171) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_283) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_283) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_287) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_287) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_273) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_273) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_164) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_164) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_171) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_171) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_283) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_283) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_375) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_375) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_407) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_407) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_164) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_164) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_171) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_171) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_417) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_417) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_287) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_287) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_407) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_407) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_164) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_164) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_171) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_171) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_463) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_463) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_287) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_287) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_273) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_273) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_164) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_164) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_171) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_171) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_287) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_287) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_184) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:117 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_184) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_512) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_512) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_535) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_535) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_539) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_539) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_543) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_543) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_547) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_547) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_551) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_551) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_535) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_535) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_558) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:285 assert (sink_ok, \"'D' channel Grant carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_558) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_539) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_539) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_566) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_566) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_570) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_570) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_547) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_547) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is denied (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:290 assert (deny_put_ok || !bundle.denied, \"'D' channel Grant is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_535) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_535) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_558) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:295 assert (sink_ok, \"'D' channel GrantData carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_558) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_539) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_539) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_566) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_566) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_570) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_570) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_603) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_603) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:300 assert (deny_get_ok || !bundle.denied, \"'D' channel GrantData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_535) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_535) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_543) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_543) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_547) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_547) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is denied (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:308 assert (deny_put_ok || !bundle.denied, \"'D' channel AccessAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_535) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_535) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_543) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_543) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_603) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_603) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:316 assert (deny_get_ok || !bundle.denied, \"'D' channel AccessAckData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_535) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_535) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_543) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_543) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_547) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_547) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is denied (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:324 assert (deny_put_ok || !bundle.denied, \"'D' channel HintAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel valid and not TL-C (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:341 assert (!bundle.b.valid, \"'B' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel valid and not TL-C (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:342 assert (!bundle.c.valid, \"'C' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel valid and not TL-C (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:343 assert (!bundle.e.valid, \"'E' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_699 & _T_703) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_699 & _T_703) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_699 & _T_707) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_699 & _T_707) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_699 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_699 & _T_711) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_699 & _T_715) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_699 & _T_715) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_699 & _T_719) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_699 & _T_719) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_748 & _T_752) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_748 & _T_752) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_748 & _T_756) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_748 & _T_756) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_748 & _T_760) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_748 & _T_760) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_748 & _T_764) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_748 & _T_764) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_748 & _T_768) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_748 & _T_768) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_748 & _T_772) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_748 & _T_772) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_817 & _T_825) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_817 & _T_825) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_832 & _T_839) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_832 & _T_839) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_846) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_846) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_859) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at ChiplinkTest.scala:221:7)\n    at Monitor.scala:479 assert (!inflight.orR || limit === UInt(0) || watchdog < limit, \"TileLink timeout expired\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_859) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLMonitor_13( 
  input         clock, 
  input         reset, 
  input         io_in_a_ready, 
  input         io_in_a_valid, 
  input  [2:0]  io_in_a_bits_opcode, 
  input  [2:0]  io_in_a_bits_param, 
  input  [2:0]  io_in_a_bits_size, 
  input  [6:0]  io_in_a_bits_source, 
  input  [28:0] io_in_a_bits_address, 
  input  [3:0]  io_in_a_bits_mask, 
  input         io_in_a_bits_corrupt, 
  input         io_in_c_ready, 
  input         io_in_c_valid, 
  input  [2:0]  io_in_c_bits_opcode, 
  input  [2:0]  io_in_c_bits_param, 
  input  [2:0]  io_in_c_bits_size, 
  input  [6:0]  io_in_c_bits_source, 
  input  [28:0] io_in_c_bits_address, 
  input         io_in_c_bits_corrupt, 
  input         io_in_d_ready, 
  input         io_in_d_valid, 
  input  [2:0]  io_in_d_bits_opcode, 
  input  [1:0]  io_in_d_bits_param, 
  input  [2:0]  io_in_d_bits_size, 
  input  [6:0]  io_in_d_bits_source, 
  input         io_in_d_bits_sink, 
  input         io_in_d_bits_denied, 
  input         io_in_d_bits_corrupt, 
  input         io_in_e_valid 
);
  wire [31:0] plusarg_reader_out; 
  wire [2:0] _T_7; 
  wire  _T_8; 
  wire  _T_16; 
  wire  _T_24; 
  wire  _T_32; 
  wire  _T_40; 
  wire  _T_48; 
  wire  _T_56; 
  wire  _T_64; 
  wire  _T_70; 
  wire  _T_71; 
  wire  _T_72; 
  wire  _T_73; 
  wire  _T_74; 
  wire  _T_75; 
  wire  _T_76; 
  wire [12:0] _T_78; 
  wire [5:0] _T_79; 
  wire [5:0] _T_80; 
  wire [28:0] _GEN_33; 
  wire [28:0] _T_81; 
  wire  _T_82; 
  wire  _T_84; 
  wire [1:0] _T_85; 
  wire [1:0] _T_87; 
  wire  _T_88; 
  wire  _T_89; 
  wire  _T_90; 
  wire  _T_91; 
  wire  _T_93; 
  wire  _T_94; 
  wire  _T_96; 
  wire  _T_97; 
  wire  _T_98; 
  wire  _T_99; 
  wire  _T_100; 
  wire  _T_101; 
  wire  _T_102; 
  wire  _T_103; 
  wire  _T_104; 
  wire  _T_105; 
  wire  _T_106; 
  wire  _T_107; 
  wire  _T_108; 
  wire  _T_109; 
  wire  _T_110; 
  wire  _T_111; 
  wire  _T_112; 
  wire [3:0] _T_115; 
  wire  _T_246; 
  wire  _T_248; 
  wire [28:0] _T_251; 
  wire [29:0] _T_252; 
  wire [29:0] _T_253; 
  wire [29:0] _T_254; 
  wire  _T_255; 
  wire  _T_256; 
  wire  _T_259; 
  wire  _T_260; 
  wire  _T_329; 
  wire  _T_346; 
  wire  _T_347; 
  wire  _T_349; 
  wire  _T_350; 
  wire  _T_353; 
  wire  _T_354; 
  wire  _T_356; 
  wire  _T_357; 
  wire  _T_358; 
  wire  _T_360; 
  wire  _T_361; 
  wire [3:0] _T_362; 
  wire  _T_363; 
  wire  _T_365; 
  wire  _T_366; 
  wire  _T_367; 
  wire  _T_369; 
  wire  _T_370; 
  wire  _T_371; 
  wire  _T_487; 
  wire  _T_489; 
  wire  _T_490; 
  wire  _T_500; 
  wire  _T_521; 
  wire  _T_523; 
  wire  _T_524; 
  wire  _T_525; 
  wire  _T_527; 
  wire  _T_528; 
  wire  _T_533; 
  wire  _T_562; 
  wire [3:0] _T_587; 
  wire [3:0] _T_588; 
  wire  _T_589; 
  wire  _T_591; 
  wire  _T_592; 
  wire  _T_593; 
  wire  _T_614; 
  wire  _T_616; 
  wire  _T_617; 
  wire  _T_622; 
  wire  _T_643; 
  wire  _T_645; 
  wire  _T_646; 
  wire  _T_651; 
  wire  _T_680; 
  wire  _T_682; 
  wire  _T_683; 
  wire [2:0] _T_686; 
  wire  _T_687; 
  wire  _T_695; 
  wire  _T_703; 
  wire  _T_711; 
  wire  _T_719; 
  wire  _T_727; 
  wire  _T_735; 
  wire  _T_743; 
  wire  _T_749; 
  wire  _T_750; 
  wire  _T_751; 
  wire  _T_752; 
  wire  _T_753; 
  wire  _T_754; 
  wire  _T_755; 
  wire  _T_756; 
  wire  _T_757; 
  wire  _T_759; 
  wire  _T_760; 
  wire  _T_761; 
  wire  _T_763; 
  wire  _T_764; 
  wire  _T_765; 
  wire  _T_767; 
  wire  _T_768; 
  wire  _T_769; 
  wire  _T_771; 
  wire  _T_772; 
  wire  _T_773; 
  wire  _T_775; 
  wire  _T_776; 
  wire  _T_777; 
  wire  _T_782; 
  wire  _T_783; 
  wire  _T_788; 
  wire  _T_790; 
  wire  _T_791; 
  wire  _T_792; 
  wire  _T_794; 
  wire  _T_795; 
  wire  _T_805; 
  wire  _T_825; 
  wire  _T_827; 
  wire  _T_828; 
  wire  _T_834; 
  wire  _T_851; 
  wire  _T_869; 
  wire [2:0] _T_1394; 
  wire  _T_1395; 
  wire  _T_1403; 
  wire  _T_1411; 
  wire  _T_1419; 
  wire  _T_1427; 
  wire  _T_1435; 
  wire  _T_1443; 
  wire  _T_1451; 
  wire  _T_1457; 
  wire  _T_1458; 
  wire  _T_1459; 
  wire  _T_1460; 
  wire  _T_1461; 
  wire  _T_1462; 
  wire  _T_1463; 
  wire [12:0] _T_1465; 
  wire [5:0] _T_1466; 
  wire [5:0] _T_1467; 
  wire [28:0] _GEN_34; 
  wire [28:0] _T_1468; 
  wire  _T_1469; 
  wire [28:0] _T_1470; 
  wire [29:0] _T_1471; 
  wire [29:0] _T_1472; 
  wire [29:0] _T_1473; 
  wire  _T_1474; 
  wire  _T_1606; 
  wire  _T_1608; 
  wire  _T_1609; 
  wire  _T_1611; 
  wire  _T_1612; 
  wire  _T_1613; 
  wire  _T_1615; 
  wire  _T_1616; 
  wire  _T_1618; 
  wire  _T_1619; 
  wire  _T_1620; 
  wire  _T_1622; 
  wire  _T_1623; 
  wire  _T_1624; 
  wire  _T_1626; 
  wire  _T_1627; 
  wire  _T_1628; 
  wire  _T_1646; 
  wire  _T_1648; 
  wire  _T_1656; 
  wire  _T_1659; 
  wire  _T_1660; 
  wire  _T_1729; 
  wire  _T_1746; 
  wire  _T_1747; 
  wire  _T_1758; 
  wire  _T_1760; 
  wire  _T_1761; 
  wire  _T_1766; 
  wire  _T_1882; 
  wire  _T_1892; 
  wire  _T_1894; 
  wire  _T_1895; 
  wire  _T_1900; 
  wire  _T_1914; 
  wire  _T_1936; 
  wire [3:0] _T_1941; 
  wire  _T_1942; 
  wire  _T_1943; 
  reg [3:0] _T_1945; 
  reg [31:0] _RAND_0;
  wire [3:0] _T_1947; 
  wire  _T_1948; 
  reg [2:0] _T_1956; 
  reg [31:0] _RAND_1;
  reg [2:0] _T_1957; 
  reg [31:0] _RAND_2;
  reg [2:0] _T_1958; 
  reg [31:0] _RAND_3;
  reg [6:0] _T_1959; 
  reg [31:0] _RAND_4;
  reg [28:0] _T_1960; 
  reg [31:0] _RAND_5;
  wire  _T_1961; 
  wire  _T_1962; 
  wire  _T_1963; 
  wire  _T_1965; 
  wire  _T_1966; 
  wire  _T_1967; 
  wire  _T_1969; 
  wire  _T_1970; 
  wire  _T_1971; 
  wire  _T_1973; 
  wire  _T_1974; 
  wire  _T_1975; 
  wire  _T_1977; 
  wire  _T_1978; 
  wire  _T_1979; 
  wire  _T_1981; 
  wire  _T_1982; 
  wire  _T_1984; 
  wire  _T_1985; 
  wire [12:0] _T_1987; 
  wire [5:0] _T_1988; 
  wire [5:0] _T_1989; 
  wire [3:0] _T_1990; 
  wire  _T_1991; 
  reg [3:0] _T_1993; 
  reg [31:0] _RAND_6;
  wire [3:0] _T_1995; 
  wire  _T_1996; 
  reg [2:0] _T_2004; 
  reg [31:0] _RAND_7;
  reg [1:0] _T_2005; 
  reg [31:0] _RAND_8;
  reg [2:0] _T_2006; 
  reg [31:0] _RAND_9;
  reg [6:0] _T_2007; 
  reg [31:0] _RAND_10;
  reg  _T_2008; 
  reg [31:0] _RAND_11;
  reg  _T_2009; 
  reg [31:0] _RAND_12;
  wire  _T_2010; 
  wire  _T_2011; 
  wire  _T_2012; 
  wire  _T_2014; 
  wire  _T_2015; 
  wire  _T_2016; 
  wire  _T_2018; 
  wire  _T_2019; 
  wire  _T_2020; 
  wire  _T_2022; 
  wire  _T_2023; 
  wire  _T_2024; 
  wire  _T_2026; 
  wire  _T_2027; 
  wire  _T_2028; 
  wire  _T_2030; 
  wire  _T_2031; 
  wire  _T_2032; 
  wire  _T_2034; 
  wire  _T_2035; 
  wire  _T_2037; 
  wire  _T_2087; 
  wire [3:0] _T_2092; 
  wire  _T_2093; 
  reg [3:0] _T_2095; 
  reg [31:0] _RAND_13;
  wire [3:0] _T_2097; 
  wire  _T_2098; 
  reg [2:0] _T_2106; 
  reg [31:0] _RAND_14;
  reg [2:0] _T_2107; 
  reg [31:0] _RAND_15;
  reg [2:0] _T_2108; 
  reg [31:0] _RAND_16;
  reg [6:0] _T_2109; 
  reg [31:0] _RAND_17;
  reg [28:0] _T_2110; 
  reg [31:0] _RAND_18;
  wire  _T_2111; 
  wire  _T_2112; 
  wire  _T_2113; 
  wire  _T_2115; 
  wire  _T_2116; 
  wire  _T_2117; 
  wire  _T_2119; 
  wire  _T_2120; 
  wire  _T_2121; 
  wire  _T_2123; 
  wire  _T_2124; 
  wire  _T_2125; 
  wire  _T_2127; 
  wire  _T_2128; 
  wire  _T_2129; 
  wire  _T_2131; 
  wire  _T_2132; 
  wire  _T_2134; 
  reg [127:0] _T_2135; 
  reg [127:0] _RAND_19;
  reg [3:0] _T_2145; 
  reg [31:0] _RAND_20;
  wire [3:0] _T_2147; 
  wire  _T_2148; 
  reg [3:0] _T_2164; 
  reg [31:0] _RAND_21;
  wire [3:0] _T_2166; 
  wire  _T_2167; 
  wire  _T_2177; 
  wire [127:0] _T_2179; 
  wire [127:0] _T_2180; 
  wire  _T_2181; 
  wire  _T_2182; 
  wire  _T_2184; 
  wire  _T_2185; 
  wire [127:0] _GEN_27; 
  wire  _T_2189; 
  wire  _T_2191; 
  wire  _T_2192; 
  wire [127:0] _T_2193; 
  wire [127:0] _T_2194; 
  wire [127:0] _T_2195; 
  wire  _T_2196; 
  wire  _T_2198; 
  wire  _T_2199; 
  wire [127:0] _GEN_28; 
  wire  _T_2200; 
  wire  _T_2201; 
  wire  _T_2202; 
  wire  _T_2203; 
  wire  _T_2205; 
  wire  _T_2206; 
  wire [127:0] _T_2207; 
  wire [127:0] _T_2208; 
  wire [127:0] _T_2209; 
  reg [31:0] _T_2210; 
  reg [31:0] _RAND_22;
  wire  _T_2211; 
  wire  _T_2212; 
  wire  _T_2213; 
  wire  _T_2214; 
  wire  _T_2215; 
  wire  _T_2216; 
  wire  _T_2218; 
  wire  _T_2219; 
  wire [31:0] _T_2221; 
  wire  _T_2224; 
  reg  _T_2225; 
  reg [31:0] _RAND_23;
  reg [3:0] _T_2234; 
  reg [31:0] _RAND_24;
  wire [3:0] _T_2236; 
  wire  _T_2237; 
  wire  _T_2247; 
  wire  _T_2248; 
  wire  _T_2249; 
  wire  _T_2250; 
  wire  _T_2251; 
  wire  _T_2252; 
  wire [1:0] _T_2253; 
  wire  _T_2254; 
  wire  _T_2256; 
  wire  _T_2258; 
  wire  _T_2259; 
  wire [1:0] _GEN_31; 
  wire  _T_2245; 
  wire  _T_2265; 
  wire  _T_2269; 
  wire  _T_2270; 
  wire [1:0] _GEN_32; 
  wire  _T_2271; 
  wire  _T_2260; 
  wire  _T_2272; 
  wire  _T_2273; 
  wire  _GEN_35; 
  wire  _GEN_51; 
  wire  _GEN_69; 
  wire  _GEN_81; 
  wire  _GEN_91; 
  wire  _GEN_101; 
  wire  _GEN_111; 
  wire  _GEN_121; 
  wire  _GEN_131; 
  wire  _GEN_141; 
  wire  _GEN_153; 
  wire  _GEN_165; 
  wire  _GEN_171; 
  wire  _GEN_177; 
  wire  _GEN_183; 
  wire  _GEN_195; 
  wire  _GEN_205; 
  wire  _GEN_219; 
  wire  _GEN_231; 
  wire  _GEN_241; 
  wire  _GEN_249; 
  dual_plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0)) plusarg_reader ( 
    .out(plusarg_reader_out)
  );
  assign _T_7 = io_in_a_bits_source[6:4]; 
  assign _T_8 = _T_7 == 3'h0; 
  assign _T_16 = _T_7 == 3'h1; 
  assign _T_24 = _T_7 == 3'h2; 
  assign _T_32 = _T_7 == 3'h3; 
  assign _T_40 = _T_7 == 3'h4; 
  assign _T_48 = _T_7 == 3'h5; 
  assign _T_56 = _T_7 == 3'h6; 
  assign _T_64 = _T_7 == 3'h7; 
  assign _T_70 = _T_8 | _T_16; 
  assign _T_71 = _T_70 | _T_24; 
  assign _T_72 = _T_71 | _T_32; 
  assign _T_73 = _T_72 | _T_40; 
  assign _T_74 = _T_73 | _T_48; 
  assign _T_75 = _T_74 | _T_56; 
  assign _T_76 = _T_75 | _T_64; 
  assign _T_78 = 13'h3f << io_in_a_bits_size; 
  assign _T_79 = _T_78[5:0]; 
  assign _T_80 = ~ _T_79; 
  assign _GEN_33 = {{23'd0}, _T_80}; 
  assign _T_81 = io_in_a_bits_address & _GEN_33; 
  assign _T_82 = _T_81 == 29'h0; 
  assign _T_84 = io_in_a_bits_size[0]; 
  assign _T_85 = 2'h1 << _T_84; 
  assign _T_87 = _T_85 | 2'h1; 
  assign _T_88 = io_in_a_bits_size >= 3'h2; 
  assign _T_89 = _T_87[1]; 
  assign _T_90 = io_in_a_bits_address[1]; 
  assign _T_91 = _T_90 == 1'h0; 
  assign _T_93 = _T_89 & _T_91; 
  assign _T_94 = _T_88 | _T_93; 
  assign _T_96 = _T_89 & _T_90; 
  assign _T_97 = _T_88 | _T_96; 
  assign _T_98 = _T_87[0]; 
  assign _T_99 = io_in_a_bits_address[0]; 
  assign _T_100 = _T_99 == 1'h0; 
  assign _T_101 = _T_91 & _T_100; 
  assign _T_102 = _T_98 & _T_101; 
  assign _T_103 = _T_94 | _T_102; 
  assign _T_104 = _T_91 & _T_99; 
  assign _T_105 = _T_98 & _T_104; 
  assign _T_106 = _T_94 | _T_105; 
  assign _T_107 = _T_90 & _T_100; 
  assign _T_108 = _T_98 & _T_107; 
  assign _T_109 = _T_97 | _T_108; 
  assign _T_110 = _T_90 & _T_99; 
  assign _T_111 = _T_98 & _T_110; 
  assign _T_112 = _T_97 | _T_111; 
  assign _T_115 = {_T_112,_T_109,_T_106,_T_103}; 
  assign _T_246 = io_in_a_bits_opcode == 3'h6; 
  assign _T_248 = io_in_a_bits_size <= 3'h6; 
  assign _T_251 = io_in_a_bits_address ^ 29'h10000000; 
  assign _T_252 = {1'b0,$signed(_T_251)}; 
  assign _T_253 = $signed(_T_252) & $signed(-30'sh10000000); 
  assign _T_254 = $signed(_T_253); 
  assign _T_255 = $signed(_T_254) == $signed(30'sh0); 
  assign _T_256 = _T_248 & _T_255; 
  assign _T_259 = _T_256 | reset; 
  assign _T_260 = _T_259 == 1'h0; 
  assign _T_329 = _T_8 ? _T_248 : 1'h0; 
  assign _T_346 = _T_329 | reset; 
  assign _T_347 = _T_346 == 1'h0; 
  assign _T_349 = _T_76 | reset; 
  assign _T_350 = _T_349 == 1'h0; 
  assign _T_353 = _T_88 | reset; 
  assign _T_354 = _T_353 == 1'h0; 
  assign _T_356 = _T_82 | reset; 
  assign _T_357 = _T_356 == 1'h0; 
  assign _T_358 = io_in_a_bits_param <= 3'h2; 
  assign _T_360 = _T_358 | reset; 
  assign _T_361 = _T_360 == 1'h0; 
  assign _T_362 = ~ io_in_a_bits_mask; 
  assign _T_363 = _T_362 == 4'h0; 
  assign _T_365 = _T_363 | reset; 
  assign _T_366 = _T_365 == 1'h0; 
  assign _T_367 = io_in_a_bits_corrupt == 1'h0; 
  assign _T_369 = _T_367 | reset; 
  assign _T_370 = _T_369 == 1'h0; 
  assign _T_371 = io_in_a_bits_opcode == 3'h7; 
  assign _T_487 = io_in_a_bits_param != 3'h0; 
  assign _T_489 = _T_487 | reset; 
  assign _T_490 = _T_489 == 1'h0; 
  assign _T_500 = io_in_a_bits_opcode == 3'h4; 
  assign _T_521 = io_in_a_bits_param == 3'h0; 
  assign _T_523 = _T_521 | reset; 
  assign _T_524 = _T_523 == 1'h0; 
  assign _T_525 = io_in_a_bits_mask == _T_115; 
  assign _T_527 = _T_525 | reset; 
  assign _T_528 = _T_527 == 1'h0; 
  assign _T_533 = io_in_a_bits_opcode == 3'h0; 
  assign _T_562 = io_in_a_bits_opcode == 3'h1; 
  assign _T_587 = ~ _T_115; 
  assign _T_588 = io_in_a_bits_mask & _T_587; 
  assign _T_589 = _T_588 == 4'h0; 
  assign _T_591 = _T_589 | reset; 
  assign _T_592 = _T_591 == 1'h0; 
  assign _T_593 = io_in_a_bits_opcode == 3'h2; 
  assign _T_614 = io_in_a_bits_param <= 3'h4; 
  assign _T_616 = _T_614 | reset; 
  assign _T_617 = _T_616 == 1'h0; 
  assign _T_622 = io_in_a_bits_opcode == 3'h3; 
  assign _T_643 = io_in_a_bits_param <= 3'h3; 
  assign _T_645 = _T_643 | reset; 
  assign _T_646 = _T_645 == 1'h0; 
  assign _T_651 = io_in_a_bits_opcode == 3'h5; 
  assign _T_680 = io_in_d_bits_opcode <= 3'h6; 
  assign _T_682 = _T_680 | reset; 
  assign _T_683 = _T_682 == 1'h0; 
  assign _T_686 = io_in_d_bits_source[6:4]; 
  assign _T_687 = _T_686 == 3'h0; 
  assign _T_695 = _T_686 == 3'h1; 
  assign _T_703 = _T_686 == 3'h2; 
  assign _T_711 = _T_686 == 3'h3; 
  assign _T_719 = _T_686 == 3'h4; 
  assign _T_727 = _T_686 == 3'h5; 
  assign _T_735 = _T_686 == 3'h6; 
  assign _T_743 = _T_686 == 3'h7; 
  assign _T_749 = _T_687 | _T_695; 
  assign _T_750 = _T_749 | _T_703; 
  assign _T_751 = _T_750 | _T_711; 
  assign _T_752 = _T_751 | _T_719; 
  assign _T_753 = _T_752 | _T_727; 
  assign _T_754 = _T_753 | _T_735; 
  assign _T_755 = _T_754 | _T_743; 
  assign _T_756 = io_in_d_bits_sink < 1'h1; 
  assign _T_757 = io_in_d_bits_opcode == 3'h6; 
  assign _T_759 = _T_755 | reset; 
  assign _T_760 = _T_759 == 1'h0; 
  assign _T_761 = io_in_d_bits_size >= 3'h2; 
  assign _T_763 = _T_761 | reset; 
  assign _T_764 = _T_763 == 1'h0; 
  assign _T_765 = io_in_d_bits_param == 2'h0; 
  assign _T_767 = _T_765 | reset; 
  assign _T_768 = _T_767 == 1'h0; 
  assign _T_769 = io_in_d_bits_corrupt == 1'h0; 
  assign _T_771 = _T_769 | reset; 
  assign _T_772 = _T_771 == 1'h0; 
  assign _T_773 = io_in_d_bits_denied == 1'h0; 
  assign _T_775 = _T_773 | reset; 
  assign _T_776 = _T_775 == 1'h0; 
  assign _T_777 = io_in_d_bits_opcode == 3'h4; 
  assign _T_782 = _T_756 | reset; 
  assign _T_783 = _T_782 == 1'h0; 
  assign _T_788 = io_in_d_bits_param <= 2'h2; 
  assign _T_790 = _T_788 | reset; 
  assign _T_791 = _T_790 == 1'h0; 
  assign _T_792 = io_in_d_bits_param != 2'h2; 
  assign _T_794 = _T_792 | reset; 
  assign _T_795 = _T_794 == 1'h0; 
  assign _T_805 = io_in_d_bits_opcode == 3'h5; 
  assign _T_825 = _T_773 | io_in_d_bits_corrupt; 
  assign _T_827 = _T_825 | reset; 
  assign _T_828 = _T_827 == 1'h0; 
  assign _T_834 = io_in_d_bits_opcode == 3'h0; 
  assign _T_851 = io_in_d_bits_opcode == 3'h1; 
  assign _T_869 = io_in_d_bits_opcode == 3'h2; 
  assign _T_1394 = io_in_c_bits_source[6:4]; 
  assign _T_1395 = _T_1394 == 3'h0; 
  assign _T_1403 = _T_1394 == 3'h1; 
  assign _T_1411 = _T_1394 == 3'h2; 
  assign _T_1419 = _T_1394 == 3'h3; 
  assign _T_1427 = _T_1394 == 3'h4; 
  assign _T_1435 = _T_1394 == 3'h5; 
  assign _T_1443 = _T_1394 == 3'h6; 
  assign _T_1451 = _T_1394 == 3'h7; 
  assign _T_1457 = _T_1395 | _T_1403; 
  assign _T_1458 = _T_1457 | _T_1411; 
  assign _T_1459 = _T_1458 | _T_1419; 
  assign _T_1460 = _T_1459 | _T_1427; 
  assign _T_1461 = _T_1460 | _T_1435; 
  assign _T_1462 = _T_1461 | _T_1443; 
  assign _T_1463 = _T_1462 | _T_1451; 
  assign _T_1465 = 13'h3f << io_in_c_bits_size; 
  assign _T_1466 = _T_1465[5:0]; 
  assign _T_1467 = ~ _T_1466; 
  assign _GEN_34 = {{23'd0}, _T_1467}; 
  assign _T_1468 = io_in_c_bits_address & _GEN_34; 
  assign _T_1469 = _T_1468 == 29'h0; 
  assign _T_1470 = io_in_c_bits_address ^ 29'h10000000; 
  assign _T_1471 = {1'b0,$signed(_T_1470)}; 
  assign _T_1472 = $signed(_T_1471) & $signed(-30'sh10000000); 
  assign _T_1473 = $signed(_T_1472); 
  assign _T_1474 = $signed(_T_1473) == $signed(30'sh0); 
  assign _T_1606 = io_in_c_bits_opcode == 3'h4; 
  assign _T_1608 = _T_1474 | reset; 
  assign _T_1609 = _T_1608 == 1'h0; 
  assign _T_1611 = _T_1463 | reset; 
  assign _T_1612 = _T_1611 == 1'h0; 
  assign _T_1613 = io_in_c_bits_size >= 3'h2; 
  assign _T_1615 = _T_1613 | reset; 
  assign _T_1616 = _T_1615 == 1'h0; 
  assign _T_1618 = _T_1469 | reset; 
  assign _T_1619 = _T_1618 == 1'h0; 
  assign _T_1620 = io_in_c_bits_param <= 3'h5; 
  assign _T_1622 = _T_1620 | reset; 
  assign _T_1623 = _T_1622 == 1'h0; 
  assign _T_1624 = io_in_c_bits_corrupt == 1'h0; 
  assign _T_1626 = _T_1624 | reset; 
  assign _T_1627 = _T_1626 == 1'h0; 
  assign _T_1628 = io_in_c_bits_opcode == 3'h5; 
  assign _T_1646 = io_in_c_bits_opcode == 3'h6; 
  assign _T_1648 = io_in_c_bits_size <= 3'h6; 
  assign _T_1656 = _T_1648 & _T_1474; 
  assign _T_1659 = _T_1656 | reset; 
  assign _T_1660 = _T_1659 == 1'h0; 
  assign _T_1729 = _T_1395 ? _T_1648 : 1'h0; 
  assign _T_1746 = _T_1729 | reset; 
  assign _T_1747 = _T_1746 == 1'h0; 
  assign _T_1758 = io_in_c_bits_param <= 3'h2; 
  assign _T_1760 = _T_1758 | reset; 
  assign _T_1761 = _T_1760 == 1'h0; 
  assign _T_1766 = io_in_c_bits_opcode == 3'h7; 
  assign _T_1882 = io_in_c_bits_opcode == 3'h0; 
  assign _T_1892 = io_in_c_bits_param == 3'h0; 
  assign _T_1894 = _T_1892 | reset; 
  assign _T_1895 = _T_1894 == 1'h0; 
  assign _T_1900 = io_in_c_bits_opcode == 3'h1; 
  assign _T_1914 = io_in_c_bits_opcode == 3'h2; 
  assign _T_1936 = io_in_a_ready & io_in_a_valid; 
  assign _T_1941 = _T_80[5:2]; 
  assign _T_1942 = io_in_a_bits_opcode[2]; 
  assign _T_1943 = _T_1942 == 1'h0; 
  assign _T_1947 = _T_1945 - 4'h1; 
  assign _T_1948 = _T_1945 == 4'h0; 
  assign _T_1961 = _T_1948 == 1'h0; 
  assign _T_1962 = io_in_a_valid & _T_1961; 
  assign _T_1963 = io_in_a_bits_opcode == _T_1956; 
  assign _T_1965 = _T_1963 | reset; 
  assign _T_1966 = _T_1965 == 1'h0; 
  assign _T_1967 = io_in_a_bits_param == _T_1957; 
  assign _T_1969 = _T_1967 | reset; 
  assign _T_1970 = _T_1969 == 1'h0; 
  assign _T_1971 = io_in_a_bits_size == _T_1958; 
  assign _T_1973 = _T_1971 | reset; 
  assign _T_1974 = _T_1973 == 1'h0; 
  assign _T_1975 = io_in_a_bits_source == _T_1959; 
  assign _T_1977 = _T_1975 | reset; 
  assign _T_1978 = _T_1977 == 1'h0; 
  assign _T_1979 = io_in_a_bits_address == _T_1960; 
  assign _T_1981 = _T_1979 | reset; 
  assign _T_1982 = _T_1981 == 1'h0; 
  assign _T_1984 = _T_1936 & _T_1948; 
  assign _T_1985 = io_in_d_ready & io_in_d_valid; 
  assign _T_1987 = 13'h3f << io_in_d_bits_size; 
  assign _T_1988 = _T_1987[5:0]; 
  assign _T_1989 = ~ _T_1988; 
  assign _T_1990 = _T_1989[5:2]; 
  assign _T_1991 = io_in_d_bits_opcode[0]; 
  assign _T_1995 = _T_1993 - 4'h1; 
  assign _T_1996 = _T_1993 == 4'h0; 
  assign _T_2010 = _T_1996 == 1'h0; 
  assign _T_2011 = io_in_d_valid & _T_2010; 
  assign _T_2012 = io_in_d_bits_opcode == _T_2004; 
  assign _T_2014 = _T_2012 | reset; 
  assign _T_2015 = _T_2014 == 1'h0; 
  assign _T_2016 = io_in_d_bits_param == _T_2005; 
  assign _T_2018 = _T_2016 | reset; 
  assign _T_2019 = _T_2018 == 1'h0; 
  assign _T_2020 = io_in_d_bits_size == _T_2006; 
  assign _T_2022 = _T_2020 | reset; 
  assign _T_2023 = _T_2022 == 1'h0; 
  assign _T_2024 = io_in_d_bits_source == _T_2007; 
  assign _T_2026 = _T_2024 | reset; 
  assign _T_2027 = _T_2026 == 1'h0; 
  assign _T_2028 = io_in_d_bits_sink == _T_2008; 
  assign _T_2030 = _T_2028 | reset; 
  assign _T_2031 = _T_2030 == 1'h0; 
  assign _T_2032 = io_in_d_bits_denied == _T_2009; 
  assign _T_2034 = _T_2032 | reset; 
  assign _T_2035 = _T_2034 == 1'h0; 
  assign _T_2037 = _T_1985 & _T_1996; 
  assign _T_2087 = io_in_c_ready & io_in_c_valid; 
  assign _T_2092 = _T_1467[5:2]; 
  assign _T_2093 = io_in_c_bits_opcode[0]; 
  assign _T_2097 = _T_2095 - 4'h1; 
  assign _T_2098 = _T_2095 == 4'h0; 
  assign _T_2111 = _T_2098 == 1'h0; 
  assign _T_2112 = io_in_c_valid & _T_2111; 
  assign _T_2113 = io_in_c_bits_opcode == _T_2106; 
  assign _T_2115 = _T_2113 | reset; 
  assign _T_2116 = _T_2115 == 1'h0; 
  assign _T_2117 = io_in_c_bits_param == _T_2107; 
  assign _T_2119 = _T_2117 | reset; 
  assign _T_2120 = _T_2119 == 1'h0; 
  assign _T_2121 = io_in_c_bits_size == _T_2108; 
  assign _T_2123 = _T_2121 | reset; 
  assign _T_2124 = _T_2123 == 1'h0; 
  assign _T_2125 = io_in_c_bits_source == _T_2109; 
  assign _T_2127 = _T_2125 | reset; 
  assign _T_2128 = _T_2127 == 1'h0; 
  assign _T_2129 = io_in_c_bits_address == _T_2110; 
  assign _T_2131 = _T_2129 | reset; 
  assign _T_2132 = _T_2131 == 1'h0; 
  assign _T_2134 = _T_2087 & _T_2098; 
  assign _T_2147 = _T_2145 - 4'h1; 
  assign _T_2148 = _T_2145 == 4'h0; 
  assign _T_2166 = _T_2164 - 4'h1; 
  assign _T_2167 = _T_2164 == 4'h0; 
  assign _T_2177 = _T_1936 & _T_2148; 
  assign _T_2179 = 128'h1 << io_in_a_bits_source; 
  assign _T_2180 = _T_2135 >> io_in_a_bits_source; 
  assign _T_2181 = _T_2180[0]; 
  assign _T_2182 = _T_2181 == 1'h0; 
  assign _T_2184 = _T_2182 | reset; 
  assign _T_2185 = _T_2184 == 1'h0; 
  assign _GEN_27 = _T_2177 ? _T_2179 : 128'h0; 
  assign _T_2189 = _T_1985 & _T_2167; 
  assign _T_2191 = _T_757 == 1'h0; 
  assign _T_2192 = _T_2189 & _T_2191; 
  assign _T_2193 = 128'h1 << io_in_d_bits_source; 
  assign _T_2194 = _GEN_27 | _T_2135; 
  assign _T_2195 = _T_2194 >> io_in_d_bits_source; 
  assign _T_2196 = _T_2195[0]; 
  assign _T_2198 = _T_2196 | reset; 
  assign _T_2199 = _T_2198 == 1'h0; 
  assign _GEN_28 = _T_2192 ? _T_2193 : 128'h0; 
  assign _T_2200 = _GEN_27 != _GEN_28; 
  assign _T_2201 = _GEN_27 != 128'h0; 
  assign _T_2202 = _T_2201 == 1'h0; 
  assign _T_2203 = _T_2200 | _T_2202; 
  assign _T_2205 = _T_2203 | reset; 
  assign _T_2206 = _T_2205 == 1'h0; 
  assign _T_2207 = _T_2135 | _GEN_27; 
  assign _T_2208 = ~ _GEN_28; 
  assign _T_2209 = _T_2207 & _T_2208; 
  assign _T_2211 = _T_2135 != 128'h0; 
  assign _T_2212 = _T_2211 == 1'h0; 
  assign _T_2213 = plusarg_reader_out == 32'h0; 
  assign _T_2214 = _T_2212 | _T_2213; 
  assign _T_2215 = _T_2210 < plusarg_reader_out; 
  assign _T_2216 = _T_2214 | _T_2215; 
  assign _T_2218 = _T_2216 | reset; 
  assign _T_2219 = _T_2218 == 1'h0; 
  assign _T_2221 = _T_2210 + 32'h1; 
  assign _T_2224 = _T_1936 | _T_1985; 
  assign _T_2236 = _T_2234 - 4'h1; 
  assign _T_2237 = _T_2234 == 4'h0; 
  assign _T_2247 = _T_1985 & _T_2237; 
  assign _T_2248 = io_in_d_bits_opcode[2]; 
  assign _T_2249 = io_in_d_bits_opcode[1]; 
  assign _T_2250 = _T_2249 == 1'h0; 
  assign _T_2251 = _T_2248 & _T_2250; 
  assign _T_2252 = _T_2247 & _T_2251; 
  assign _T_2253 = 2'h1 << io_in_d_bits_sink; 
  assign _T_2254 = _T_2225 >> io_in_d_bits_sink; 
  assign _T_2256 = _T_2254 == 1'h0; 
  assign _T_2258 = _T_2256 | reset; 
  assign _T_2259 = _T_2258 == 1'h0; 
  assign _GEN_31 = _T_2252 ? _T_2253 : 2'h0; 
  assign _T_2245 = _GEN_31[0]; 
  assign _T_2265 = _T_2245 | _T_2225; 
  assign _T_2269 = _T_2265 | reset; 
  assign _T_2270 = _T_2269 == 1'h0; 
  assign _GEN_32 = io_in_e_valid ? 2'h1 : 2'h0; 
  assign _T_2271 = _T_2225 | _T_2245; 
  assign _T_2260 = _GEN_32[0]; 
  assign _T_2272 = ~ _T_2260; 
  assign _T_2273 = _T_2271 & _T_2272; 
  assign _GEN_35 = io_in_a_valid & _T_246; 
  assign _GEN_51 = io_in_a_valid & _T_371; 
  assign _GEN_69 = io_in_a_valid & _T_500; 
  assign _GEN_81 = io_in_a_valid & _T_533; 
  assign _GEN_91 = io_in_a_valid & _T_562; 
  assign _GEN_101 = io_in_a_valid & _T_593; 
  assign _GEN_111 = io_in_a_valid & _T_622; 
  assign _GEN_121 = io_in_a_valid & _T_651; 
  assign _GEN_131 = io_in_d_valid & _T_757; 
  assign _GEN_141 = io_in_d_valid & _T_777; 
  assign _GEN_153 = io_in_d_valid & _T_805; 
  assign _GEN_165 = io_in_d_valid & _T_834; 
  assign _GEN_171 = io_in_d_valid & _T_851; 
  assign _GEN_177 = io_in_d_valid & _T_869; 
  assign _GEN_183 = io_in_c_valid & _T_1606; 
  assign _GEN_195 = io_in_c_valid & _T_1628; 
  assign _GEN_205 = io_in_c_valid & _T_1646; 
  assign _GEN_219 = io_in_c_valid & _T_1766; 
  assign _GEN_231 = io_in_c_valid & _T_1882; 
  assign _GEN_241 = io_in_c_valid & _T_1900; 
  assign _GEN_249 = io_in_c_valid & _T_1914; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1945 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1956 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1957 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1958 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1959 = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1960 = _RAND_5[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_1993 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_2004 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_2005 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_2006 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_2007 = _RAND_10[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_2008 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_2009 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_2095 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_2106 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_2107 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_2108 = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_2109 = _RAND_17[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_2110 = _RAND_18[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {4{`RANDOM}};
  _T_2135 = _RAND_19[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_2145 = _RAND_20[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_2164 = _RAND_21[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_2210 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_2225 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_2234 = _RAND_24[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_1945 <= 4'h0;
    end else begin
      if (_T_1936) begin
        if (_T_1948) begin
          if (_T_1943) begin
            _T_1945 <= _T_1941;
          end else begin
            _T_1945 <= 4'h0;
          end
        end else begin
          _T_1945 <= _T_1947;
        end
      end
    end
    if (_T_1984) begin
      _T_1956 <= io_in_a_bits_opcode;
    end
    if (_T_1984) begin
      _T_1957 <= io_in_a_bits_param;
    end
    if (_T_1984) begin
      _T_1958 <= io_in_a_bits_size;
    end
    if (_T_1984) begin
      _T_1959 <= io_in_a_bits_source;
    end
    if (_T_1984) begin
      _T_1960 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_1993 <= 4'h0;
    end else begin
      if (_T_1985) begin
        if (_T_1996) begin
          if (_T_1991) begin
            _T_1993 <= _T_1990;
          end else begin
            _T_1993 <= 4'h0;
          end
        end else begin
          _T_1993 <= _T_1995;
        end
      end
    end
    if (_T_2037) begin
      _T_2004 <= io_in_d_bits_opcode;
    end
    if (_T_2037) begin
      _T_2005 <= io_in_d_bits_param;
    end
    if (_T_2037) begin
      _T_2006 <= io_in_d_bits_size;
    end
    if (_T_2037) begin
      _T_2007 <= io_in_d_bits_source;
    end
    if (_T_2037) begin
      _T_2008 <= io_in_d_bits_sink;
    end
    if (_T_2037) begin
      _T_2009 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_2095 <= 4'h0;
    end else begin
      if (_T_2087) begin
        if (_T_2098) begin
          if (_T_2093) begin
            _T_2095 <= _T_2092;
          end else begin
            _T_2095 <= 4'h0;
          end
        end else begin
          _T_2095 <= _T_2097;
        end
      end
    end
    if (_T_2134) begin
      _T_2106 <= io_in_c_bits_opcode;
    end
    if (_T_2134) begin
      _T_2107 <= io_in_c_bits_param;
    end
    if (_T_2134) begin
      _T_2108 <= io_in_c_bits_size;
    end
    if (_T_2134) begin
      _T_2109 <= io_in_c_bits_source;
    end
    if (_T_2134) begin
      _T_2110 <= io_in_c_bits_address;
    end
    if (reset) begin
      _T_2135 <= 128'h0;
    end else begin
      _T_2135 <= _T_2209;
    end
    if (reset) begin
      _T_2145 <= 4'h0;
    end else begin
      if (_T_1936) begin
        if (_T_2148) begin
          if (_T_1943) begin
            _T_2145 <= _T_1941;
          end else begin
            _T_2145 <= 4'h0;
          end
        end else begin
          _T_2145 <= _T_2147;
        end
      end
    end
    if (reset) begin
      _T_2164 <= 4'h0;
    end else begin
      if (_T_1985) begin
        if (_T_2167) begin
          if (_T_1991) begin
            _T_2164 <= _T_1990;
          end else begin
            _T_2164 <= 4'h0;
          end
        end else begin
          _T_2164 <= _T_2166;
        end
      end
    end
    if (reset) begin
      _T_2210 <= 32'h0;
    end else begin
      if (_T_2224) begin
        _T_2210 <= 32'h0;
      end else begin
        _T_2210 <= _T_2221;
      end
    end
    if (reset) begin
      _T_2225 <= 1'h0;
    end else begin
      _T_2225 <= _T_2273;
    end
    if (reset) begin
      _T_2234 <= 4'h0;
    end else begin
      if (_T_1985) begin
        if (_T_2237) begin
          if (_T_1991) begin
            _T_2234 <= _T_1990;
          end else begin
            _T_2234 <= 4'h0;
          end
        end else begin
          _T_2234 <= _T_2236;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel has invalid opcode (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:39 assert (TLMessages.isA(bundle.opcode), \"'A' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:46 assert (visible(edge.address(bundle), bundle.source, edge), \"'A' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_260) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_260) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_347) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_347) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_350) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_350) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_354) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_354) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_357) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_357) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_361) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_361) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_366) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_366) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_370) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:56 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_370) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_260) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_260) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_347) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_347) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_350) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_350) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_354) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_354) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_357) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_357) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_361) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_361) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_490) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_490) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_366) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_366) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_370) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:68 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_370) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_260) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & _T_260) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_350) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & _T_350) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_357) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & _T_357) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_524) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & _T_524) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_528) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & _T_528) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_370) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:77 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & _T_370) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_81 & _T_260) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_81 & _T_260) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_81 & _T_350) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_81 & _T_350) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_81 & _T_357) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_81 & _T_357) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_81 & _T_524) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_81 & _T_524) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_81 & _T_528) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_81 & _T_528) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_260) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_260) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_350) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_350) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_357) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_357) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_524) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_524) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_592) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_592) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_260) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_260) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_350) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_350) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_357) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_357) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_617) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_617) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_528) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_528) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & _T_260) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & _T_260) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & _T_350) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & _T_350) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & _T_357) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & _T_357) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & _T_646) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & _T_646) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & _T_528) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & _T_528) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_260) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_260) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_350) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_350) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_357) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_357) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_528) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_528) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_370) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:117 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_370) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_683) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_683) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_760) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_760) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_764) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_764) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_768) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_768) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_772) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_772) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_776) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_776) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_760) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_760) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_783) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:285 assert (sink_ok, \"'D' channel Grant carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_783) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_764) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_764) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_791) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_791) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_795) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_795) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_772) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_772) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is denied (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:290 assert (deny_put_ok || !bundle.denied, \"'D' channel Grant is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_760) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_760) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_783) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:295 assert (sink_ok, \"'D' channel GrantData carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_783) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_764) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_764) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_791) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_791) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_795) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_795) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_828) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_828) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:300 assert (deny_get_ok || !bundle.denied, \"'D' channel GrantData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & _T_760) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & _T_760) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & _T_768) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & _T_768) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & _T_772) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & _T_772) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is denied (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:308 assert (deny_put_ok || !bundle.denied, \"'D' channel AccessAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_760) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_760) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_768) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_768) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_828) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_828) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:316 assert (deny_get_ok || !bundle.denied, \"'D' channel AccessAckData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_177 & _T_760) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_177 & _T_760) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_177 & _T_768) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_177 & _T_768) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_177 & _T_772) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_177 & _T_772) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is denied (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:324 assert (deny_put_ok || !bundle.denied, \"'D' channel HintAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel has invalid opcode (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:122 assert (TLMessages.isB(bundle.opcode), \"'B' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:124 assert (visible(edge.address(bundle), bundle.source, edge), \"'B' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Probe type unsupported by client (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:133 assert (edge.client.supportsProbe(bundle.source, bundle.size), \"'B' channel carries Probe type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:134 assert (address_ok, \"'B' channel Probe carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries source that is not first source (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:135 assert (legal_source, \"'B' channel Probe carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:136 assert (is_aligned, \"'B' channel Probe address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:137 assert (TLPermissions.isCap(bundle.param), \"'B' channel Probe carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe contains invalid mask (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:138 assert (bundle.mask === mask, \"'B' channel Probe contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe is corrupt (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:139 assert (!bundle.corrupt, \"'B' channel Probe is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Get type unsupported by client (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:143 assert (edge.client.supportsGet(bundle.source, bundle.size), \"'B' channel carries Get type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries unmanaged address (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:144 assert (address_ok, \"'B' channel Get carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries source that is not first source (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:145 assert (legal_source, \"'B' channel Get carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:146 assert (is_aligned, \"'B' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries invalid param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:147 assert (bundle.param === UInt(0), \"'B' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get contains invalid mask (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:148 assert (bundle.mask === mask, \"'B' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get is corrupt (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:149 assert (!bundle.corrupt, \"'B' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutFull type unsupported by client (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:153 assert (edge.client.supportsPutFull(bundle.source, bundle.size), \"'B' channel carries PutFull type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries unmanaged address (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:154 assert (address_ok, \"'B' channel PutFull carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries source that is not first source (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:155 assert (legal_source, \"'B' channel PutFull carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:156 assert (is_aligned, \"'B' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries invalid param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:157 assert (bundle.param === UInt(0), \"'B' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull contains invalid mask (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:158 assert (bundle.mask === mask, \"'B' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutPartial type unsupported by client (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:162 assert (edge.client.supportsPutPartial(bundle.source, bundle.size), \"'B' channel carries PutPartial type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:163 assert (address_ok, \"'B' channel PutPartial carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:164 assert (legal_source, \"'B' channel PutPartial carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:165 assert (is_aligned, \"'B' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries invalid param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:166 assert (bundle.param === UInt(0), \"'B' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial contains invalid mask (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:167 assert ((bundle.mask & ~mask) === UInt(0), \"'B' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Arithmetic type unsupported by client (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:171 assert (edge.client.supportsArithmetic(bundle.source, bundle.size), \"'B' channel carries Arithmetic type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:172 assert (address_ok, \"'B' channel Arithmetic carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:173 assert (legal_source, \"'B' channel Arithmetic carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:174 assert (is_aligned, \"'B' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries invalid opcode param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:175 assert (TLAtomics.isArithmetic(bundle.param), \"'B' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:176 assert (bundle.mask === mask, \"'B' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Logical type unsupported by client (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:180 assert (edge.client.supportsLogical(bundle.source, bundle.size), \"'B' channel carries Logical type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries unmanaged address (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:181 assert (address_ok, \"'B' channel Logical carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries source that is not first source (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:182 assert (legal_source, \"'B' channel Logical carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:183 assert (is_aligned, \"'B' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries invalid opcode param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:184 assert (TLAtomics.isLogical(bundle.param), \"'B' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical contains invalid mask (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:185 assert (bundle.mask === mask, \"'B' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Hint type unsupported by client (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:189 assert (edge.client.supportsHint(bundle.source, bundle.size), \"'B' channel carries Hint type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries unmanaged address (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:190 assert (address_ok, \"'B' channel Hint carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries source that is not first source (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:191 assert (legal_source, \"'B' channel Hint carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:192 assert (is_aligned, \"'B' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint contains invalid mask (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:193 assert (bundle.mask === mask, \"'B' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint is corrupt (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:194 assert (!bundle.corrupt, \"'B' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel has invalid opcode (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:199 assert (TLMessages.isC(bundle.opcode), \"'C' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:205 assert (visible(edge.address(bundle), bundle.source, edge), \"'C' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_1609) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:208 assert (address_ok, \"'C' channel ProbeAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_1609) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_1612) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:209 assert (source_ok, \"'C' channel ProbeAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_1612) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_1616) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:210 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_1616) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_1619) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:211 assert (is_aligned, \"'C' channel ProbeAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_1619) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_1623) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:212 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAck carries invalid report param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_1623) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_1627) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck is corrupt (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:213 assert (!bundle.corrupt, \"'C' channel ProbeAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_1627) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1609) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:217 assert (address_ok, \"'C' channel ProbeAckData carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1609) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1612) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:218 assert (source_ok, \"'C' channel ProbeAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1612) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1616) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:219 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAckData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1616) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1619) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:220 assert (is_aligned, \"'C' channel ProbeAckData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1619) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1623) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:221 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAckData carries invalid report param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1623) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1660) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:225 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries Release type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1660) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1747) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:226 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1747) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1612) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:227 assert (source_ok, \"'C' channel Release carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1612) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1616) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:228 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel Release smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1616) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1619) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:229 assert (is_aligned, \"'C' channel Release address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1619) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1761) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid shrink param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:230 assert (TLPermissions.isShrink(bundle.param), \"'C' channel Release carries invalid shrink param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1761) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1627) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release is corrupt (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:231 assert (!bundle.corrupt, \"'C' channel Release is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1627) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1660) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:235 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries ReleaseData type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1660) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1747) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:236 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1747) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1612) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:237 assert (source_ok, \"'C' channel ReleaseData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1612) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1616) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:238 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ReleaseData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1616) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1619) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:239 assert (is_aligned, \"'C' channel ReleaseData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1619) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1761) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid shrink param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:240 assert (TLPermissions.isShrink(bundle.param), \"'C' channel ReleaseData carries invalid shrink param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1761) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1609) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:244 assert (address_ok, \"'C' channel AccessAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1609) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1612) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:245 assert (source_ok, \"'C' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1612) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1619) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:246 assert (is_aligned, \"'C' channel AccessAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1619) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1895) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:247 assert (bundle.param === UInt(0), \"'C' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1895) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1627) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck is corrupt (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:248 assert (!bundle.corrupt, \"'C' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1627) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1609) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:252 assert (address_ok, \"'C' channel AccessAckData carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1609) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1612) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:253 assert (source_ok, \"'C' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1612) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1619) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:254 assert (is_aligned, \"'C' channel AccessAckData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1619) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1895) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:255 assert (bundle.param === UInt(0), \"'C' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1895) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_249 & _T_1609) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:259 assert (address_ok, \"'C' channel HintAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_249 & _T_1609) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_249 & _T_1612) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:260 assert (source_ok, \"'C' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_249 & _T_1612) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_249 & _T_1619) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:261 assert (is_aligned, \"'C' channel HintAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_249 & _T_1619) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_249 & _T_1895) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:262 assert (bundle.param === UInt(0), \"'C' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_249 & _T_1895) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_249 & _T_1627) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck is corrupt (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:263 assert (!bundle.corrupt, \"'C' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_249 & _T_1627) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channels carries invalid sink ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:330 assert (sink_ok, \"'E' channels carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1962 & _T_1966) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1962 & _T_1966) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1962 & _T_1970) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1962 & _T_1970) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1962 & _T_1974) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1962 & _T_1974) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1962 & _T_1978) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1962 & _T_1978) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1962 & _T_1982) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1962 & _T_1982) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2011 & _T_2015) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2011 & _T_2015) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2011 & _T_2019) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2011 & _T_2019) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2011 & _T_2023) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2011 & _T_2023) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2011 & _T_2027) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2011 & _T_2027) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2011 & _T_2031) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2011 & _T_2031) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2011 & _T_2035) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2011 & _T_2035) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:378 assert (b.bits.opcode === opcode, \"'B' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:379 assert (b.bits.param  === param,  \"'B' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel size changed within multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:380 assert (b.bits.size   === size,   \"'B' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel source changed within multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:381 assert (b.bits.source === source, \"'B' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:382 assert (b.bits.address=== address,\"'B' channel addresss changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2112 & _T_2116) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:401 assert (c.bits.opcode === opcode, \"'C' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2112 & _T_2116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2112 & _T_2120) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:402 assert (c.bits.param  === param,  \"'C' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2112 & _T_2120) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2112 & _T_2124) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:403 assert (c.bits.size   === size,   \"'C' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2112 & _T_2124) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2112 & _T_2128) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:404 assert (c.bits.source === source, \"'C' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2112 & _T_2128) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2112 & _T_2132) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:405 assert (c.bits.address=== address,\"'C' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2112 & _T_2132) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2177 & _T_2185) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2177 & _T_2185) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2192 & _T_2199) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2192 & _T_2199) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2206) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2206) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2219) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:479 assert (!inflight.orR || limit === UInt(0) || watchdog < limit, \"TileLink timeout expired\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2219) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2252 & _T_2259) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:494 assert(!inflight(bundle.d.bits.sink), \"'D' channel re-used a sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2252 & _T_2259) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_e_valid & _T_2270) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at ChiplinkTest.scala:363:12)\n    at Monitor.scala:500 assert((d_set | inflight)(bundle.e.bits.sink), \"'E' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_e_valid & _T_2270) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLMonitor_14( 
  input         clock, 
  input         reset, 
  input         io_in_a_ready, 
  input         io_in_a_valid, 
  input  [2:0]  io_in_a_bits_opcode, 
  input  [2:0]  io_in_a_bits_param, 
  input  [3:0]  io_in_a_bits_size, 
  input  [6:0]  io_in_a_bits_source, 
  input  [31:0] io_in_a_bits_address, 
  input  [7:0]  io_in_a_bits_mask, 
  input         io_in_c_ready, 
  input         io_in_c_valid, 
  input  [2:0]  io_in_c_bits_opcode, 
  input  [2:0]  io_in_c_bits_param, 
  input  [3:0]  io_in_c_bits_size, 
  input  [6:0]  io_in_c_bits_source, 
  input  [31:0] io_in_c_bits_address, 
  input         io_in_c_bits_corrupt, 
  input         io_in_d_ready, 
  input         io_in_d_valid, 
  input  [2:0]  io_in_d_bits_opcode, 
  input  [1:0]  io_in_d_bits_param, 
  input  [3:0]  io_in_d_bits_size, 
  input  [6:0]  io_in_d_bits_source, 
  input         io_in_d_bits_sink, 
  input         io_in_d_bits_denied, 
  input         io_in_d_bits_corrupt, 
  input         io_in_e_ready, 
  input         io_in_e_valid, 
  input         io_in_e_bits_sink 
);
  wire [31:0] plusarg_reader_out; 
  wire [2:0] _T_7; 
  wire  _T_8; 
  wire  _T_16; 
  wire  _T_24; 
  wire  _T_32; 
  wire  _T_40; 
  wire  _T_48; 
  wire  _T_56; 
  wire  _T_64; 
  wire  _T_70; 
  wire  _T_71; 
  wire  _T_72; 
  wire  _T_73; 
  wire  _T_74; 
  wire  _T_75; 
  wire  _T_76; 
  wire [22:0] _T_78; 
  wire [7:0] _T_79; 
  wire [7:0] _T_80; 
  wire [31:0] _GEN_33; 
  wire [31:0] _T_81; 
  wire  _T_82; 
  wire [1:0] _T_84; 
  wire [3:0] _T_85; 
  wire [2:0] _T_86; 
  wire [2:0] _T_87; 
  wire  _T_88; 
  wire  _T_89; 
  wire  _T_90; 
  wire  _T_91; 
  wire  _T_93; 
  wire  _T_94; 
  wire  _T_96; 
  wire  _T_97; 
  wire  _T_98; 
  wire  _T_99; 
  wire  _T_100; 
  wire  _T_101; 
  wire  _T_102; 
  wire  _T_103; 
  wire  _T_104; 
  wire  _T_105; 
  wire  _T_106; 
  wire  _T_107; 
  wire  _T_108; 
  wire  _T_109; 
  wire  _T_110; 
  wire  _T_111; 
  wire  _T_112; 
  wire  _T_113; 
  wire  _T_114; 
  wire  _T_115; 
  wire  _T_116; 
  wire  _T_117; 
  wire  _T_118; 
  wire  _T_119; 
  wire  _T_120; 
  wire  _T_121; 
  wire  _T_122; 
  wire  _T_123; 
  wire  _T_124; 
  wire  _T_125; 
  wire  _T_126; 
  wire  _T_127; 
  wire  _T_128; 
  wire  _T_129; 
  wire  _T_130; 
  wire  _T_131; 
  wire  _T_132; 
  wire  _T_133; 
  wire  _T_134; 
  wire  _T_135; 
  wire  _T_136; 
  wire  _T_137; 
  wire  _T_138; 
  wire  _T_139; 
  wire [7:0] _T_146; 
  wire  _T_277; 
  wire [31:0] _T_279; 
  wire [32:0] _T_280; 
  wire [32:0] _T_281; 
  wire [32:0] _T_282; 
  wire  _T_283; 
  wire [31:0] _T_284; 
  wire [32:0] _T_285; 
  wire [32:0] _T_286; 
  wire [32:0] _T_287; 
  wire  _T_288; 
  wire  _T_289; 
  wire  _T_292; 
  wire [31:0] _T_295; 
  wire [32:0] _T_296; 
  wire [32:0] _T_297; 
  wire [32:0] _T_298; 
  wire  _T_299; 
  wire  _T_300; 
  wire  _T_304; 
  wire  _T_305; 
  wire  _T_374; 
  wire  _T_391; 
  wire  _T_392; 
  wire  _T_394; 
  wire  _T_395; 
  wire  _T_398; 
  wire  _T_399; 
  wire  _T_401; 
  wire  _T_402; 
  wire  _T_403; 
  wire  _T_405; 
  wire  _T_406; 
  wire [7:0] _T_407; 
  wire  _T_408; 
  wire  _T_410; 
  wire  _T_411; 
  wire  _T_416; 
  wire  _T_546; 
  wire  _T_548; 
  wire  _T_549; 
  wire  _T_559; 
  wire  _T_580; 
  wire  _T_581; 
  wire  _T_584; 
  wire  _T_585; 
  wire  _T_592; 
  wire  _T_594; 
  wire  _T_595; 
  wire  _T_596; 
  wire  _T_598; 
  wire  _T_599; 
  wire  _T_604; 
  wire  _T_619; 
  wire  _T_620; 
  wire  _T_622; 
  wire  _T_630; 
  wire  _T_632; 
  wire  _T_634; 
  wire  _T_635; 
  wire  _T_650; 
  wire [7:0] _T_692; 
  wire [7:0] _T_693; 
  wire  _T_694; 
  wire  _T_696; 
  wire  _T_697; 
  wire  _T_698; 
  wire  _T_700; 
  wire  _T_720; 
  wire  _T_723; 
  wire  _T_724; 
  wire  _T_731; 
  wire  _T_733; 
  wire  _T_734; 
  wire  _T_739; 
  wire  _T_772; 
  wire  _T_774; 
  wire  _T_775; 
  wire  _T_780; 
  wire  _T_823; 
  wire  _T_825; 
  wire  _T_826; 
  wire [2:0] _T_829; 
  wire  _T_830; 
  wire  _T_838; 
  wire  _T_846; 
  wire  _T_854; 
  wire  _T_862; 
  wire  _T_870; 
  wire  _T_878; 
  wire  _T_886; 
  wire  _T_892; 
  wire  _T_893; 
  wire  _T_894; 
  wire  _T_895; 
  wire  _T_896; 
  wire  _T_897; 
  wire  _T_898; 
  wire  _T_899; 
  wire  _T_900; 
  wire  _T_902; 
  wire  _T_903; 
  wire  _T_904; 
  wire  _T_906; 
  wire  _T_907; 
  wire  _T_908; 
  wire  _T_910; 
  wire  _T_911; 
  wire  _T_912; 
  wire  _T_914; 
  wire  _T_915; 
  wire  _T_916; 
  wire  _T_918; 
  wire  _T_919; 
  wire  _T_920; 
  wire  _T_925; 
  wire  _T_926; 
  wire  _T_931; 
  wire  _T_933; 
  wire  _T_934; 
  wire  _T_935; 
  wire  _T_937; 
  wire  _T_938; 
  wire  _T_948; 
  wire  _T_968; 
  wire  _T_970; 
  wire  _T_971; 
  wire  _T_977; 
  wire  _T_994; 
  wire  _T_1012; 
  wire [2:0] _T_1580; 
  wire  _T_1581; 
  wire  _T_1589; 
  wire  _T_1597; 
  wire  _T_1605; 
  wire  _T_1613; 
  wire  _T_1621; 
  wire  _T_1629; 
  wire  _T_1637; 
  wire  _T_1643; 
  wire  _T_1644; 
  wire  _T_1645; 
  wire  _T_1646; 
  wire  _T_1647; 
  wire  _T_1648; 
  wire  _T_1649; 
  wire [22:0] _T_1651; 
  wire [7:0] _T_1652; 
  wire [7:0] _T_1653; 
  wire [31:0] _GEN_34; 
  wire [31:0] _T_1654; 
  wire  _T_1655; 
  wire [31:0] _T_1656; 
  wire [32:0] _T_1657; 
  wire [32:0] _T_1658; 
  wire [32:0] _T_1659; 
  wire  _T_1660; 
  wire [31:0] _T_1661; 
  wire [32:0] _T_1662; 
  wire [32:0] _T_1663; 
  wire [32:0] _T_1664; 
  wire  _T_1665; 
  wire [31:0] _T_1666; 
  wire [32:0] _T_1667; 
  wire [32:0] _T_1668; 
  wire [32:0] _T_1669; 
  wire  _T_1670; 
  wire  _T_1672; 
  wire  _T_1673; 
  wire  _T_1804; 
  wire  _T_1806; 
  wire  _T_1807; 
  wire  _T_1809; 
  wire  _T_1810; 
  wire  _T_1811; 
  wire  _T_1813; 
  wire  _T_1814; 
  wire  _T_1816; 
  wire  _T_1817; 
  wire  _T_1818; 
  wire  _T_1820; 
  wire  _T_1821; 
  wire  _T_1822; 
  wire  _T_1824; 
  wire  _T_1825; 
  wire  _T_1826; 
  wire  _T_1844; 
  wire  _T_1859; 
  wire  _T_1867; 
  wire  _T_1871; 
  wire  _T_1872; 
  wire  _T_1941; 
  wire  _T_1958; 
  wire  _T_1959; 
  wire  _T_1970; 
  wire  _T_1972; 
  wire  _T_1973; 
  wire  _T_1978; 
  wire  _T_2108; 
  wire  _T_2118; 
  wire  _T_2120; 
  wire  _T_2121; 
  wire  _T_2126; 
  wire  _T_2140; 
  wire  _T_2158; 
  wire  _T_2160; 
  wire  _T_2161; 
  wire  _T_2162; 
  wire [4:0] _T_2167; 
  wire  _T_2168; 
  wire  _T_2169; 
  reg [4:0] _T_2171; 
  reg [31:0] _RAND_0;
  wire [4:0] _T_2173; 
  wire  _T_2174; 
  reg [2:0] _T_2182; 
  reg [31:0] _RAND_1;
  reg [2:0] _T_2183; 
  reg [31:0] _RAND_2;
  reg [3:0] _T_2184; 
  reg [31:0] _RAND_3;
  reg [6:0] _T_2185; 
  reg [31:0] _RAND_4;
  reg [31:0] _T_2186; 
  reg [31:0] _RAND_5;
  wire  _T_2187; 
  wire  _T_2188; 
  wire  _T_2189; 
  wire  _T_2191; 
  wire  _T_2192; 
  wire  _T_2193; 
  wire  _T_2195; 
  wire  _T_2196; 
  wire  _T_2197; 
  wire  _T_2199; 
  wire  _T_2200; 
  wire  _T_2201; 
  wire  _T_2203; 
  wire  _T_2204; 
  wire  _T_2205; 
  wire  _T_2207; 
  wire  _T_2208; 
  wire  _T_2210; 
  wire  _T_2211; 
  wire [22:0] _T_2213; 
  wire [7:0] _T_2214; 
  wire [7:0] _T_2215; 
  wire [4:0] _T_2216; 
  wire  _T_2217; 
  reg [4:0] _T_2219; 
  reg [31:0] _RAND_6;
  wire [4:0] _T_2221; 
  wire  _T_2222; 
  reg [2:0] _T_2230; 
  reg [31:0] _RAND_7;
  reg [1:0] _T_2231; 
  reg [31:0] _RAND_8;
  reg [3:0] _T_2232; 
  reg [31:0] _RAND_9;
  reg [6:0] _T_2233; 
  reg [31:0] _RAND_10;
  reg  _T_2234; 
  reg [31:0] _RAND_11;
  reg  _T_2235; 
  reg [31:0] _RAND_12;
  wire  _T_2236; 
  wire  _T_2237; 
  wire  _T_2238; 
  wire  _T_2240; 
  wire  _T_2241; 
  wire  _T_2242; 
  wire  _T_2244; 
  wire  _T_2245; 
  wire  _T_2246; 
  wire  _T_2248; 
  wire  _T_2249; 
  wire  _T_2250; 
  wire  _T_2252; 
  wire  _T_2253; 
  wire  _T_2254; 
  wire  _T_2256; 
  wire  _T_2257; 
  wire  _T_2258; 
  wire  _T_2260; 
  wire  _T_2261; 
  wire  _T_2263; 
  wire  _T_2313; 
  wire [4:0] _T_2318; 
  wire  _T_2319; 
  reg [4:0] _T_2321; 
  reg [31:0] _RAND_13;
  wire [4:0] _T_2323; 
  wire  _T_2324; 
  reg [2:0] _T_2332; 
  reg [31:0] _RAND_14;
  reg [2:0] _T_2333; 
  reg [31:0] _RAND_15;
  reg [3:0] _T_2334; 
  reg [31:0] _RAND_16;
  reg [6:0] _T_2335; 
  reg [31:0] _RAND_17;
  reg [31:0] _T_2336; 
  reg [31:0] _RAND_18;
  wire  _T_2337; 
  wire  _T_2338; 
  wire  _T_2339; 
  wire  _T_2341; 
  wire  _T_2342; 
  wire  _T_2343; 
  wire  _T_2345; 
  wire  _T_2346; 
  wire  _T_2347; 
  wire  _T_2349; 
  wire  _T_2350; 
  wire  _T_2351; 
  wire  _T_2353; 
  wire  _T_2354; 
  wire  _T_2355; 
  wire  _T_2357; 
  wire  _T_2358; 
  wire  _T_2360; 
  reg [127:0] _T_2361; 
  reg [127:0] _RAND_19;
  reg [4:0] _T_2371; 
  reg [31:0] _RAND_20;
  wire [4:0] _T_2373; 
  wire  _T_2374; 
  reg [4:0] _T_2390; 
  reg [31:0] _RAND_21;
  wire [4:0] _T_2392; 
  wire  _T_2393; 
  wire  _T_2403; 
  wire [127:0] _T_2405; 
  wire [127:0] _T_2406; 
  wire  _T_2407; 
  wire  _T_2408; 
  wire  _T_2410; 
  wire  _T_2411; 
  wire [127:0] _GEN_27; 
  wire  _T_2415; 
  wire  _T_2417; 
  wire  _T_2418; 
  wire [127:0] _T_2419; 
  wire [127:0] _T_2420; 
  wire [127:0] _T_2421; 
  wire  _T_2422; 
  wire  _T_2424; 
  wire  _T_2425; 
  wire [127:0] _GEN_28; 
  wire  _T_2426; 
  wire  _T_2427; 
  wire  _T_2428; 
  wire  _T_2429; 
  wire  _T_2431; 
  wire  _T_2432; 
  wire [127:0] _T_2433; 
  wire [127:0] _T_2434; 
  wire [127:0] _T_2435; 
  reg [31:0] _T_2436; 
  reg [31:0] _RAND_22;
  wire  _T_2437; 
  wire  _T_2438; 
  wire  _T_2439; 
  wire  _T_2440; 
  wire  _T_2441; 
  wire  _T_2442; 
  wire  _T_2444; 
  wire  _T_2445; 
  wire [31:0] _T_2447; 
  wire  _T_2450; 
  reg  _T_2451; 
  reg [31:0] _RAND_23;
  reg [4:0] _T_2460; 
  reg [31:0] _RAND_24;
  wire [4:0] _T_2462; 
  wire  _T_2463; 
  wire  _T_2473; 
  wire  _T_2474; 
  wire  _T_2475; 
  wire  _T_2476; 
  wire  _T_2477; 
  wire  _T_2478; 
  wire [1:0] _T_2479; 
  wire  _T_2480; 
  wire  _T_2482; 
  wire  _T_2484; 
  wire  _T_2485; 
  wire [1:0] _GEN_31; 
  wire  _T_2487; 
  wire [1:0] _T_2490; 
  wire  _T_2471; 
  wire  _T_2491; 
  wire  _T_2492; 
  wire  _T_2495; 
  wire  _T_2496; 
  wire [1:0] _GEN_32; 
  wire  _T_2497; 
  wire  _T_2486; 
  wire  _T_2498; 
  wire  _T_2499; 
  wire  _GEN_35; 
  wire  _GEN_49; 
  wire  _GEN_65; 
  wire  _GEN_75; 
  wire  _GEN_85; 
  wire  _GEN_95; 
  wire  _GEN_105; 
  wire  _GEN_115; 
  wire  _GEN_123; 
  wire  _GEN_133; 
  wire  _GEN_145; 
  wire  _GEN_157; 
  wire  _GEN_163; 
  wire  _GEN_169; 
  wire  _GEN_175; 
  wire  _GEN_187; 
  wire  _GEN_197; 
  wire  _GEN_211; 
  wire  _GEN_223; 
  wire  _GEN_233; 
  wire  _GEN_241; 
  dual_plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0)) plusarg_reader ( 
    .out(plusarg_reader_out)
  );
  assign _T_7 = io_in_a_bits_source[6:4]; 
  assign _T_8 = _T_7 == 3'h0; 
  assign _T_16 = _T_7 == 3'h1; 
  assign _T_24 = _T_7 == 3'h2; 
  assign _T_32 = _T_7 == 3'h3; 
  assign _T_40 = _T_7 == 3'h4; 
  assign _T_48 = _T_7 == 3'h5; 
  assign _T_56 = _T_7 == 3'h6; 
  assign _T_64 = _T_7 == 3'h7; 
  assign _T_70 = _T_8 | _T_16; 
  assign _T_71 = _T_70 | _T_24; 
  assign _T_72 = _T_71 | _T_32; 
  assign _T_73 = _T_72 | _T_40; 
  assign _T_74 = _T_73 | _T_48; 
  assign _T_75 = _T_74 | _T_56; 
  assign _T_76 = _T_75 | _T_64; 
  assign _T_78 = 23'hff << io_in_a_bits_size; 
  assign _T_79 = _T_78[7:0]; 
  assign _T_80 = ~ _T_79; 
  assign _GEN_33 = {{24'd0}, _T_80}; 
  assign _T_81 = io_in_a_bits_address & _GEN_33; 
  assign _T_82 = _T_81 == 32'h0; 
  assign _T_84 = io_in_a_bits_size[1:0]; 
  assign _T_85 = 4'h1 << _T_84; 
  assign _T_86 = _T_85[2:0]; 
  assign _T_87 = _T_86 | 3'h1; 
  assign _T_88 = io_in_a_bits_size >= 4'h3; 
  assign _T_89 = _T_87[2]; 
  assign _T_90 = io_in_a_bits_address[2]; 
  assign _T_91 = _T_90 == 1'h0; 
  assign _T_93 = _T_89 & _T_91; 
  assign _T_94 = _T_88 | _T_93; 
  assign _T_96 = _T_89 & _T_90; 
  assign _T_97 = _T_88 | _T_96; 
  assign _T_98 = _T_87[1]; 
  assign _T_99 = io_in_a_bits_address[1]; 
  assign _T_100 = _T_99 == 1'h0; 
  assign _T_101 = _T_91 & _T_100; 
  assign _T_102 = _T_98 & _T_101; 
  assign _T_103 = _T_94 | _T_102; 
  assign _T_104 = _T_91 & _T_99; 
  assign _T_105 = _T_98 & _T_104; 
  assign _T_106 = _T_94 | _T_105; 
  assign _T_107 = _T_90 & _T_100; 
  assign _T_108 = _T_98 & _T_107; 
  assign _T_109 = _T_97 | _T_108; 
  assign _T_110 = _T_90 & _T_99; 
  assign _T_111 = _T_98 & _T_110; 
  assign _T_112 = _T_97 | _T_111; 
  assign _T_113 = _T_87[0]; 
  assign _T_114 = io_in_a_bits_address[0]; 
  assign _T_115 = _T_114 == 1'h0; 
  assign _T_116 = _T_101 & _T_115; 
  assign _T_117 = _T_113 & _T_116; 
  assign _T_118 = _T_103 | _T_117; 
  assign _T_119 = _T_101 & _T_114; 
  assign _T_120 = _T_113 & _T_119; 
  assign _T_121 = _T_103 | _T_120; 
  assign _T_122 = _T_104 & _T_115; 
  assign _T_123 = _T_113 & _T_122; 
  assign _T_124 = _T_106 | _T_123; 
  assign _T_125 = _T_104 & _T_114; 
  assign _T_126 = _T_113 & _T_125; 
  assign _T_127 = _T_106 | _T_126; 
  assign _T_128 = _T_107 & _T_115; 
  assign _T_129 = _T_113 & _T_128; 
  assign _T_130 = _T_109 | _T_129; 
  assign _T_131 = _T_107 & _T_114; 
  assign _T_132 = _T_113 & _T_131; 
  assign _T_133 = _T_109 | _T_132; 
  assign _T_134 = _T_110 & _T_115; 
  assign _T_135 = _T_113 & _T_134; 
  assign _T_136 = _T_112 | _T_135; 
  assign _T_137 = _T_110 & _T_114; 
  assign _T_138 = _T_113 & _T_137; 
  assign _T_139 = _T_112 | _T_138; 
  assign _T_146 = {_T_139,_T_136,_T_133,_T_130,_T_127,_T_124,_T_121,_T_118}; 
  assign _T_277 = io_in_a_bits_opcode == 3'h6; 
  assign _T_279 = io_in_a_bits_address ^ 32'h80000000; 
  assign _T_280 = {1'b0,$signed(_T_279)}; 
  assign _T_281 = $signed(_T_280) & $signed(-33'sh80000000); 
  assign _T_282 = $signed(_T_281); 
  assign _T_283 = $signed(_T_282) == $signed(33'sh0); 
  assign _T_284 = io_in_a_bits_address ^ 32'h40000000; 
  assign _T_285 = {1'b0,$signed(_T_284)}; 
  assign _T_286 = $signed(_T_285) & $signed(-33'sh20000000); 
  assign _T_287 = $signed(_T_286); 
  assign _T_288 = $signed(_T_287) == $signed(33'sh0); 
  assign _T_289 = _T_283 | _T_288; 
  assign _T_292 = io_in_a_bits_size <= 4'h6; 
  assign _T_295 = io_in_a_bits_address ^ 32'h10000000; 
  assign _T_296 = {1'b0,$signed(_T_295)}; 
  assign _T_297 = $signed(_T_296) & $signed(-33'sh10000000); 
  assign _T_298 = $signed(_T_297); 
  assign _T_299 = $signed(_T_298) == $signed(33'sh0); 
  assign _T_300 = _T_292 & _T_299; 
  assign _T_304 = _T_300 | reset; 
  assign _T_305 = _T_304 == 1'h0; 
  assign _T_374 = _T_8 ? _T_292 : 1'h0; 
  assign _T_391 = _T_374 | reset; 
  assign _T_392 = _T_391 == 1'h0; 
  assign _T_394 = _T_76 | reset; 
  assign _T_395 = _T_394 == 1'h0; 
  assign _T_398 = _T_88 | reset; 
  assign _T_399 = _T_398 == 1'h0; 
  assign _T_401 = _T_82 | reset; 
  assign _T_402 = _T_401 == 1'h0; 
  assign _T_403 = io_in_a_bits_param <= 3'h2; 
  assign _T_405 = _T_403 | reset; 
  assign _T_406 = _T_405 == 1'h0; 
  assign _T_407 = ~ io_in_a_bits_mask; 
  assign _T_408 = _T_407 == 8'h0; 
  assign _T_410 = _T_408 | reset; 
  assign _T_411 = _T_410 == 1'h0; 
  assign _T_416 = io_in_a_bits_opcode == 3'h7; 
  assign _T_546 = io_in_a_bits_param != 3'h0; 
  assign _T_548 = _T_546 | reset; 
  assign _T_549 = _T_548 == 1'h0; 
  assign _T_559 = io_in_a_bits_opcode == 3'h4; 
  assign _T_580 = _T_289 | _T_299; 
  assign _T_581 = _T_292 & _T_580; 
  assign _T_584 = _T_581 | reset; 
  assign _T_585 = _T_584 == 1'h0; 
  assign _T_592 = io_in_a_bits_param == 3'h0; 
  assign _T_594 = _T_592 | reset; 
  assign _T_595 = _T_594 == 1'h0; 
  assign _T_596 = io_in_a_bits_mask == _T_146; 
  assign _T_598 = _T_596 | reset; 
  assign _T_599 = _T_598 == 1'h0; 
  assign _T_604 = io_in_a_bits_opcode == 3'h0; 
  assign _T_619 = _T_283 | _T_299; 
  assign _T_620 = _T_292 & _T_619; 
  assign _T_622 = io_in_a_bits_size <= 4'h8; 
  assign _T_630 = _T_622 & _T_288; 
  assign _T_632 = _T_620 | _T_630; 
  assign _T_634 = _T_632 | reset; 
  assign _T_635 = _T_634 == 1'h0; 
  assign _T_650 = io_in_a_bits_opcode == 3'h1; 
  assign _T_692 = ~ _T_146; 
  assign _T_693 = io_in_a_bits_mask & _T_692; 
  assign _T_694 = _T_693 == 8'h0; 
  assign _T_696 = _T_694 | reset; 
  assign _T_697 = _T_696 == 1'h0; 
  assign _T_698 = io_in_a_bits_opcode == 3'h2; 
  assign _T_700 = io_in_a_bits_size <= 4'h3; 
  assign _T_720 = _T_700 & _T_580; 
  assign _T_723 = _T_720 | reset; 
  assign _T_724 = _T_723 == 1'h0; 
  assign _T_731 = io_in_a_bits_param <= 3'h4; 
  assign _T_733 = _T_731 | reset; 
  assign _T_734 = _T_733 == 1'h0; 
  assign _T_739 = io_in_a_bits_opcode == 3'h3; 
  assign _T_772 = io_in_a_bits_param <= 3'h3; 
  assign _T_774 = _T_772 | reset; 
  assign _T_775 = _T_774 == 1'h0; 
  assign _T_780 = io_in_a_bits_opcode == 3'h5; 
  assign _T_823 = io_in_d_bits_opcode <= 3'h6; 
  assign _T_825 = _T_823 | reset; 
  assign _T_826 = _T_825 == 1'h0; 
  assign _T_829 = io_in_d_bits_source[6:4]; 
  assign _T_830 = _T_829 == 3'h0; 
  assign _T_838 = _T_829 == 3'h1; 
  assign _T_846 = _T_829 == 3'h2; 
  assign _T_854 = _T_829 == 3'h3; 
  assign _T_862 = _T_829 == 3'h4; 
  assign _T_870 = _T_829 == 3'h5; 
  assign _T_878 = _T_829 == 3'h6; 
  assign _T_886 = _T_829 == 3'h7; 
  assign _T_892 = _T_830 | _T_838; 
  assign _T_893 = _T_892 | _T_846; 
  assign _T_894 = _T_893 | _T_854; 
  assign _T_895 = _T_894 | _T_862; 
  assign _T_896 = _T_895 | _T_870; 
  assign _T_897 = _T_896 | _T_878; 
  assign _T_898 = _T_897 | _T_886; 
  assign _T_899 = io_in_d_bits_sink < 1'h1; 
  assign _T_900 = io_in_d_bits_opcode == 3'h6; 
  assign _T_902 = _T_898 | reset; 
  assign _T_903 = _T_902 == 1'h0; 
  assign _T_904 = io_in_d_bits_size >= 4'h3; 
  assign _T_906 = _T_904 | reset; 
  assign _T_907 = _T_906 == 1'h0; 
  assign _T_908 = io_in_d_bits_param == 2'h0; 
  assign _T_910 = _T_908 | reset; 
  assign _T_911 = _T_910 == 1'h0; 
  assign _T_912 = io_in_d_bits_corrupt == 1'h0; 
  assign _T_914 = _T_912 | reset; 
  assign _T_915 = _T_914 == 1'h0; 
  assign _T_916 = io_in_d_bits_denied == 1'h0; 
  assign _T_918 = _T_916 | reset; 
  assign _T_919 = _T_918 == 1'h0; 
  assign _T_920 = io_in_d_bits_opcode == 3'h4; 
  assign _T_925 = _T_899 | reset; 
  assign _T_926 = _T_925 == 1'h0; 
  assign _T_931 = io_in_d_bits_param <= 2'h2; 
  assign _T_933 = _T_931 | reset; 
  assign _T_934 = _T_933 == 1'h0; 
  assign _T_935 = io_in_d_bits_param != 2'h2; 
  assign _T_937 = _T_935 | reset; 
  assign _T_938 = _T_937 == 1'h0; 
  assign _T_948 = io_in_d_bits_opcode == 3'h5; 
  assign _T_968 = _T_916 | io_in_d_bits_corrupt; 
  assign _T_970 = _T_968 | reset; 
  assign _T_971 = _T_970 == 1'h0; 
  assign _T_977 = io_in_d_bits_opcode == 3'h0; 
  assign _T_994 = io_in_d_bits_opcode == 3'h1; 
  assign _T_1012 = io_in_d_bits_opcode == 3'h2; 
  assign _T_1580 = io_in_c_bits_source[6:4]; 
  assign _T_1581 = _T_1580 == 3'h0; 
  assign _T_1589 = _T_1580 == 3'h1; 
  assign _T_1597 = _T_1580 == 3'h2; 
  assign _T_1605 = _T_1580 == 3'h3; 
  assign _T_1613 = _T_1580 == 3'h4; 
  assign _T_1621 = _T_1580 == 3'h5; 
  assign _T_1629 = _T_1580 == 3'h6; 
  assign _T_1637 = _T_1580 == 3'h7; 
  assign _T_1643 = _T_1581 | _T_1589; 
  assign _T_1644 = _T_1643 | _T_1597; 
  assign _T_1645 = _T_1644 | _T_1605; 
  assign _T_1646 = _T_1645 | _T_1613; 
  assign _T_1647 = _T_1646 | _T_1621; 
  assign _T_1648 = _T_1647 | _T_1629; 
  assign _T_1649 = _T_1648 | _T_1637; 
  assign _T_1651 = 23'hff << io_in_c_bits_size; 
  assign _T_1652 = _T_1651[7:0]; 
  assign _T_1653 = ~ _T_1652; 
  assign _GEN_34 = {{24'd0}, _T_1653}; 
  assign _T_1654 = io_in_c_bits_address & _GEN_34; 
  assign _T_1655 = _T_1654 == 32'h0; 
  assign _T_1656 = io_in_c_bits_address ^ 32'h80000000; 
  assign _T_1657 = {1'b0,$signed(_T_1656)}; 
  assign _T_1658 = $signed(_T_1657) & $signed(-33'sh80000000); 
  assign _T_1659 = $signed(_T_1658); 
  assign _T_1660 = $signed(_T_1659) == $signed(33'sh0); 
  assign _T_1661 = io_in_c_bits_address ^ 32'h40000000; 
  assign _T_1662 = {1'b0,$signed(_T_1661)}; 
  assign _T_1663 = $signed(_T_1662) & $signed(-33'sh20000000); 
  assign _T_1664 = $signed(_T_1663); 
  assign _T_1665 = $signed(_T_1664) == $signed(33'sh0); 
  assign _T_1666 = io_in_c_bits_address ^ 32'h10000000; 
  assign _T_1667 = {1'b0,$signed(_T_1666)}; 
  assign _T_1668 = $signed(_T_1667) & $signed(-33'sh10000000); 
  assign _T_1669 = $signed(_T_1668); 
  assign _T_1670 = $signed(_T_1669) == $signed(33'sh0); 
  assign _T_1672 = _T_1660 | _T_1665; 
  assign _T_1673 = _T_1672 | _T_1670; 
  assign _T_1804 = io_in_c_bits_opcode == 3'h4; 
  assign _T_1806 = _T_1673 | reset; 
  assign _T_1807 = _T_1806 == 1'h0; 
  assign _T_1809 = _T_1649 | reset; 
  assign _T_1810 = _T_1809 == 1'h0; 
  assign _T_1811 = io_in_c_bits_size >= 4'h3; 
  assign _T_1813 = _T_1811 | reset; 
  assign _T_1814 = _T_1813 == 1'h0; 
  assign _T_1816 = _T_1655 | reset; 
  assign _T_1817 = _T_1816 == 1'h0; 
  assign _T_1818 = io_in_c_bits_param <= 3'h5; 
  assign _T_1820 = _T_1818 | reset; 
  assign _T_1821 = _T_1820 == 1'h0; 
  assign _T_1822 = io_in_c_bits_corrupt == 1'h0; 
  assign _T_1824 = _T_1822 | reset; 
  assign _T_1825 = _T_1824 == 1'h0; 
  assign _T_1826 = io_in_c_bits_opcode == 3'h5; 
  assign _T_1844 = io_in_c_bits_opcode == 3'h6; 
  assign _T_1859 = io_in_c_bits_size <= 4'h6; 
  assign _T_1867 = _T_1859 & _T_1670; 
  assign _T_1871 = _T_1867 | reset; 
  assign _T_1872 = _T_1871 == 1'h0; 
  assign _T_1941 = _T_1581 ? _T_1859 : 1'h0; 
  assign _T_1958 = _T_1941 | reset; 
  assign _T_1959 = _T_1958 == 1'h0; 
  assign _T_1970 = io_in_c_bits_param <= 3'h2; 
  assign _T_1972 = _T_1970 | reset; 
  assign _T_1973 = _T_1972 == 1'h0; 
  assign _T_1978 = io_in_c_bits_opcode == 3'h7; 
  assign _T_2108 = io_in_c_bits_opcode == 3'h0; 
  assign _T_2118 = io_in_c_bits_param == 3'h0; 
  assign _T_2120 = _T_2118 | reset; 
  assign _T_2121 = _T_2120 == 1'h0; 
  assign _T_2126 = io_in_c_bits_opcode == 3'h1; 
  assign _T_2140 = io_in_c_bits_opcode == 3'h2; 
  assign _T_2158 = io_in_e_bits_sink < 1'h1; 
  assign _T_2160 = _T_2158 | reset; 
  assign _T_2161 = _T_2160 == 1'h0; 
  assign _T_2162 = io_in_a_ready & io_in_a_valid; 
  assign _T_2167 = _T_80[7:3]; 
  assign _T_2168 = io_in_a_bits_opcode[2]; 
  assign _T_2169 = _T_2168 == 1'h0; 
  assign _T_2173 = _T_2171 - 5'h1; 
  assign _T_2174 = _T_2171 == 5'h0; 
  assign _T_2187 = _T_2174 == 1'h0; 
  assign _T_2188 = io_in_a_valid & _T_2187; 
  assign _T_2189 = io_in_a_bits_opcode == _T_2182; 
  assign _T_2191 = _T_2189 | reset; 
  assign _T_2192 = _T_2191 == 1'h0; 
  assign _T_2193 = io_in_a_bits_param == _T_2183; 
  assign _T_2195 = _T_2193 | reset; 
  assign _T_2196 = _T_2195 == 1'h0; 
  assign _T_2197 = io_in_a_bits_size == _T_2184; 
  assign _T_2199 = _T_2197 | reset; 
  assign _T_2200 = _T_2199 == 1'h0; 
  assign _T_2201 = io_in_a_bits_source == _T_2185; 
  assign _T_2203 = _T_2201 | reset; 
  assign _T_2204 = _T_2203 == 1'h0; 
  assign _T_2205 = io_in_a_bits_address == _T_2186; 
  assign _T_2207 = _T_2205 | reset; 
  assign _T_2208 = _T_2207 == 1'h0; 
  assign _T_2210 = _T_2162 & _T_2174; 
  assign _T_2211 = io_in_d_ready & io_in_d_valid; 
  assign _T_2213 = 23'hff << io_in_d_bits_size; 
  assign _T_2214 = _T_2213[7:0]; 
  assign _T_2215 = ~ _T_2214; 
  assign _T_2216 = _T_2215[7:3]; 
  assign _T_2217 = io_in_d_bits_opcode[0]; 
  assign _T_2221 = _T_2219 - 5'h1; 
  assign _T_2222 = _T_2219 == 5'h0; 
  assign _T_2236 = _T_2222 == 1'h0; 
  assign _T_2237 = io_in_d_valid & _T_2236; 
  assign _T_2238 = io_in_d_bits_opcode == _T_2230; 
  assign _T_2240 = _T_2238 | reset; 
  assign _T_2241 = _T_2240 == 1'h0; 
  assign _T_2242 = io_in_d_bits_param == _T_2231; 
  assign _T_2244 = _T_2242 | reset; 
  assign _T_2245 = _T_2244 == 1'h0; 
  assign _T_2246 = io_in_d_bits_size == _T_2232; 
  assign _T_2248 = _T_2246 | reset; 
  assign _T_2249 = _T_2248 == 1'h0; 
  assign _T_2250 = io_in_d_bits_source == _T_2233; 
  assign _T_2252 = _T_2250 | reset; 
  assign _T_2253 = _T_2252 == 1'h0; 
  assign _T_2254 = io_in_d_bits_sink == _T_2234; 
  assign _T_2256 = _T_2254 | reset; 
  assign _T_2257 = _T_2256 == 1'h0; 
  assign _T_2258 = io_in_d_bits_denied == _T_2235; 
  assign _T_2260 = _T_2258 | reset; 
  assign _T_2261 = _T_2260 == 1'h0; 
  assign _T_2263 = _T_2211 & _T_2222; 
  assign _T_2313 = io_in_c_ready & io_in_c_valid; 
  assign _T_2318 = _T_1653[7:3]; 
  assign _T_2319 = io_in_c_bits_opcode[0]; 
  assign _T_2323 = _T_2321 - 5'h1; 
  assign _T_2324 = _T_2321 == 5'h0; 
  assign _T_2337 = _T_2324 == 1'h0; 
  assign _T_2338 = io_in_c_valid & _T_2337; 
  assign _T_2339 = io_in_c_bits_opcode == _T_2332; 
  assign _T_2341 = _T_2339 | reset; 
  assign _T_2342 = _T_2341 == 1'h0; 
  assign _T_2343 = io_in_c_bits_param == _T_2333; 
  assign _T_2345 = _T_2343 | reset; 
  assign _T_2346 = _T_2345 == 1'h0; 
  assign _T_2347 = io_in_c_bits_size == _T_2334; 
  assign _T_2349 = _T_2347 | reset; 
  assign _T_2350 = _T_2349 == 1'h0; 
  assign _T_2351 = io_in_c_bits_source == _T_2335; 
  assign _T_2353 = _T_2351 | reset; 
  assign _T_2354 = _T_2353 == 1'h0; 
  assign _T_2355 = io_in_c_bits_address == _T_2336; 
  assign _T_2357 = _T_2355 | reset; 
  assign _T_2358 = _T_2357 == 1'h0; 
  assign _T_2360 = _T_2313 & _T_2324; 
  assign _T_2373 = _T_2371 - 5'h1; 
  assign _T_2374 = _T_2371 == 5'h0; 
  assign _T_2392 = _T_2390 - 5'h1; 
  assign _T_2393 = _T_2390 == 5'h0; 
  assign _T_2403 = _T_2162 & _T_2374; 
  assign _T_2405 = 128'h1 << io_in_a_bits_source; 
  assign _T_2406 = _T_2361 >> io_in_a_bits_source; 
  assign _T_2407 = _T_2406[0]; 
  assign _T_2408 = _T_2407 == 1'h0; 
  assign _T_2410 = _T_2408 | reset; 
  assign _T_2411 = _T_2410 == 1'h0; 
  assign _GEN_27 = _T_2403 ? _T_2405 : 128'h0; 
  assign _T_2415 = _T_2211 & _T_2393; 
  assign _T_2417 = _T_900 == 1'h0; 
  assign _T_2418 = _T_2415 & _T_2417; 
  assign _T_2419 = 128'h1 << io_in_d_bits_source; 
  assign _T_2420 = _GEN_27 | _T_2361; 
  assign _T_2421 = _T_2420 >> io_in_d_bits_source; 
  assign _T_2422 = _T_2421[0]; 
  assign _T_2424 = _T_2422 | reset; 
  assign _T_2425 = _T_2424 == 1'h0; 
  assign _GEN_28 = _T_2418 ? _T_2419 : 128'h0; 
  assign _T_2426 = _GEN_27 != _GEN_28; 
  assign _T_2427 = _GEN_27 != 128'h0; 
  assign _T_2428 = _T_2427 == 1'h0; 
  assign _T_2429 = _T_2426 | _T_2428; 
  assign _T_2431 = _T_2429 | reset; 
  assign _T_2432 = _T_2431 == 1'h0; 
  assign _T_2433 = _T_2361 | _GEN_27; 
  assign _T_2434 = ~ _GEN_28; 
  assign _T_2435 = _T_2433 & _T_2434; 
  assign _T_2437 = _T_2361 != 128'h0; 
  assign _T_2438 = _T_2437 == 1'h0; 
  assign _T_2439 = plusarg_reader_out == 32'h0; 
  assign _T_2440 = _T_2438 | _T_2439; 
  assign _T_2441 = _T_2436 < plusarg_reader_out; 
  assign _T_2442 = _T_2440 | _T_2441; 
  assign _T_2444 = _T_2442 | reset; 
  assign _T_2445 = _T_2444 == 1'h0; 
  assign _T_2447 = _T_2436 + 32'h1; 
  assign _T_2450 = _T_2162 | _T_2211; 
  assign _T_2462 = _T_2460 - 5'h1; 
  assign _T_2463 = _T_2460 == 5'h0; 
  assign _T_2473 = _T_2211 & _T_2463; 
  assign _T_2474 = io_in_d_bits_opcode[2]; 
  assign _T_2475 = io_in_d_bits_opcode[1]; 
  assign _T_2476 = _T_2475 == 1'h0; 
  assign _T_2477 = _T_2474 & _T_2476; 
  assign _T_2478 = _T_2473 & _T_2477; 
  assign _T_2479 = 2'h1 << io_in_d_bits_sink; 
  assign _T_2480 = _T_2451 >> io_in_d_bits_sink; 
  assign _T_2482 = _T_2480 == 1'h0; 
  assign _T_2484 = _T_2482 | reset; 
  assign _T_2485 = _T_2484 == 1'h0; 
  assign _GEN_31 = _T_2478 ? _T_2479 : 2'h0; 
  assign _T_2487 = io_in_e_ready & io_in_e_valid; 
  assign _T_2490 = 2'h1 << io_in_e_bits_sink; 
  assign _T_2471 = _GEN_31[0]; 
  assign _T_2491 = _T_2471 | _T_2451; 
  assign _T_2492 = _T_2491 >> io_in_e_bits_sink; 
  assign _T_2495 = _T_2492 | reset; 
  assign _T_2496 = _T_2495 == 1'h0; 
  assign _GEN_32 = _T_2487 ? _T_2490 : 2'h0; 
  assign _T_2497 = _T_2451 | _T_2471; 
  assign _T_2486 = _GEN_32[0]; 
  assign _T_2498 = ~ _T_2486; 
  assign _T_2499 = _T_2497 & _T_2498; 
  assign _GEN_35 = io_in_a_valid & _T_277; 
  assign _GEN_49 = io_in_a_valid & _T_416; 
  assign _GEN_65 = io_in_a_valid & _T_559; 
  assign _GEN_75 = io_in_a_valid & _T_604; 
  assign _GEN_85 = io_in_a_valid & _T_650; 
  assign _GEN_95 = io_in_a_valid & _T_698; 
  assign _GEN_105 = io_in_a_valid & _T_739; 
  assign _GEN_115 = io_in_a_valid & _T_780; 
  assign _GEN_123 = io_in_d_valid & _T_900; 
  assign _GEN_133 = io_in_d_valid & _T_920; 
  assign _GEN_145 = io_in_d_valid & _T_948; 
  assign _GEN_157 = io_in_d_valid & _T_977; 
  assign _GEN_163 = io_in_d_valid & _T_994; 
  assign _GEN_169 = io_in_d_valid & _T_1012; 
  assign _GEN_175 = io_in_c_valid & _T_1804; 
  assign _GEN_187 = io_in_c_valid & _T_1826; 
  assign _GEN_197 = io_in_c_valid & _T_1844; 
  assign _GEN_211 = io_in_c_valid & _T_1978; 
  assign _GEN_223 = io_in_c_valid & _T_2108; 
  assign _GEN_233 = io_in_c_valid & _T_2126; 
  assign _GEN_241 = io_in_c_valid & _T_2140; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2171 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_2182 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2183 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_2184 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_2185 = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_2186 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_2219 = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_2230 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_2231 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_2232 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_2233 = _RAND_10[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_2234 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_2235 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_2321 = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_2332 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_2333 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_2334 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_2335 = _RAND_17[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_2336 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {4{`RANDOM}};
  _T_2361 = _RAND_19[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_2371 = _RAND_20[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_2390 = _RAND_21[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_2436 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_2451 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_2460 = _RAND_24[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_2171 <= 5'h0;
    end else begin
      if (_T_2162) begin
        if (_T_2174) begin
          if (_T_2169) begin
            _T_2171 <= _T_2167;
          end else begin
            _T_2171 <= 5'h0;
          end
        end else begin
          _T_2171 <= _T_2173;
        end
      end
    end
    if (_T_2210) begin
      _T_2182 <= io_in_a_bits_opcode;
    end
    if (_T_2210) begin
      _T_2183 <= io_in_a_bits_param;
    end
    if (_T_2210) begin
      _T_2184 <= io_in_a_bits_size;
    end
    if (_T_2210) begin
      _T_2185 <= io_in_a_bits_source;
    end
    if (_T_2210) begin
      _T_2186 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_2219 <= 5'h0;
    end else begin
      if (_T_2211) begin
        if (_T_2222) begin
          if (_T_2217) begin
            _T_2219 <= _T_2216;
          end else begin
            _T_2219 <= 5'h0;
          end
        end else begin
          _T_2219 <= _T_2221;
        end
      end
    end
    if (_T_2263) begin
      _T_2230 <= io_in_d_bits_opcode;
    end
    if (_T_2263) begin
      _T_2231 <= io_in_d_bits_param;
    end
    if (_T_2263) begin
      _T_2232 <= io_in_d_bits_size;
    end
    if (_T_2263) begin
      _T_2233 <= io_in_d_bits_source;
    end
    if (_T_2263) begin
      _T_2234 <= io_in_d_bits_sink;
    end
    if (_T_2263) begin
      _T_2235 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_2321 <= 5'h0;
    end else begin
      if (_T_2313) begin
        if (_T_2324) begin
          if (_T_2319) begin
            _T_2321 <= _T_2318;
          end else begin
            _T_2321 <= 5'h0;
          end
        end else begin
          _T_2321 <= _T_2323;
        end
      end
    end
    if (_T_2360) begin
      _T_2332 <= io_in_c_bits_opcode;
    end
    if (_T_2360) begin
      _T_2333 <= io_in_c_bits_param;
    end
    if (_T_2360) begin
      _T_2334 <= io_in_c_bits_size;
    end
    if (_T_2360) begin
      _T_2335 <= io_in_c_bits_source;
    end
    if (_T_2360) begin
      _T_2336 <= io_in_c_bits_address;
    end
    if (reset) begin
      _T_2361 <= 128'h0;
    end else begin
      _T_2361 <= _T_2435;
    end
    if (reset) begin
      _T_2371 <= 5'h0;
    end else begin
      if (_T_2162) begin
        if (_T_2374) begin
          if (_T_2169) begin
            _T_2371 <= _T_2167;
          end else begin
            _T_2371 <= 5'h0;
          end
        end else begin
          _T_2371 <= _T_2373;
        end
      end
    end
    if (reset) begin
      _T_2390 <= 5'h0;
    end else begin
      if (_T_2211) begin
        if (_T_2393) begin
          if (_T_2217) begin
            _T_2390 <= _T_2216;
          end else begin
            _T_2390 <= 5'h0;
          end
        end else begin
          _T_2390 <= _T_2392;
        end
      end
    end
    if (reset) begin
      _T_2436 <= 32'h0;
    end else begin
      if (_T_2450) begin
        _T_2436 <= 32'h0;
      end else begin
        _T_2436 <= _T_2447;
      end
    end
    if (reset) begin
      _T_2451 <= 1'h0;
    end else begin
      _T_2451 <= _T_2499;
    end
    if (reset) begin
      _T_2460 <= 5'h0;
    end else begin
      if (_T_2211) begin
        if (_T_2463) begin
          if (_T_2217) begin
            _T_2460 <= _T_2216;
          end else begin
            _T_2460 <= 5'h0;
          end
        end else begin
          _T_2460 <= _T_2462;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel has invalid opcode (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:39 assert (TLMessages.isA(bundle.opcode), \"'A' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:46 assert (visible(edge.address(bundle), bundle.source, edge), \"'A' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_305) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_305) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_392) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_392) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_399) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_399) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_406) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_406) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_411) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_411) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:56 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_305) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_305) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_392) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_392) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_399) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_399) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_406) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_406) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_549) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_549) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_411) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_411) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:68 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_585) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_585) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_595) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_595) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_599) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:77 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_635) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_635) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_595) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_595) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_599) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_635) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_635) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_595) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_595) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_697) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_697) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_724) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_724) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_734) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_734) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_599) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_724) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_724) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_775) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_775) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_599) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_305) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_305) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_599) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:117 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_826) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_826) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_903) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_903) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_907) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_907) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_911) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_911) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_915) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_915) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_919) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_919) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_903) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_903) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_926) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:285 assert (sink_ok, \"'D' channel Grant carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_926) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_907) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_907) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_934) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_934) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_938) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_938) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_915) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_915) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is denied (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:290 assert (deny_put_ok || !bundle.denied, \"'D' channel Grant is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_903) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_903) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_926) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:295 assert (sink_ok, \"'D' channel GrantData carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_926) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_907) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_907) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_934) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_934) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_938) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_938) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_971) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_971) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:300 assert (deny_get_ok || !bundle.denied, \"'D' channel GrantData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_157 & _T_903) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_157 & _T_903) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_157 & _T_911) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_157 & _T_911) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_157 & _T_915) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_157 & _T_915) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is denied (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:308 assert (deny_put_ok || !bundle.denied, \"'D' channel AccessAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_903) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_903) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_911) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_911) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_971) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_971) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:316 assert (deny_get_ok || !bundle.denied, \"'D' channel AccessAckData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_169 & _T_903) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_169 & _T_903) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_169 & _T_911) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_169 & _T_911) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_169 & _T_915) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_169 & _T_915) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is denied (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:324 assert (deny_put_ok || !bundle.denied, \"'D' channel HintAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel has invalid opcode (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:122 assert (TLMessages.isB(bundle.opcode), \"'B' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:124 assert (visible(edge.address(bundle), bundle.source, edge), \"'B' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Probe type unsupported by client (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:133 assert (edge.client.supportsProbe(bundle.source, bundle.size), \"'B' channel carries Probe type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:134 assert (address_ok, \"'B' channel Probe carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries source that is not first source (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:135 assert (legal_source, \"'B' channel Probe carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:136 assert (is_aligned, \"'B' channel Probe address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:137 assert (TLPermissions.isCap(bundle.param), \"'B' channel Probe carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe contains invalid mask (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:138 assert (bundle.mask === mask, \"'B' channel Probe contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe is corrupt (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:139 assert (!bundle.corrupt, \"'B' channel Probe is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Get type unsupported by client (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:143 assert (edge.client.supportsGet(bundle.source, bundle.size), \"'B' channel carries Get type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries unmanaged address (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:144 assert (address_ok, \"'B' channel Get carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries source that is not first source (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:145 assert (legal_source, \"'B' channel Get carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:146 assert (is_aligned, \"'B' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries invalid param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:147 assert (bundle.param === UInt(0), \"'B' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get contains invalid mask (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:148 assert (bundle.mask === mask, \"'B' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get is corrupt (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:149 assert (!bundle.corrupt, \"'B' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutFull type unsupported by client (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:153 assert (edge.client.supportsPutFull(bundle.source, bundle.size), \"'B' channel carries PutFull type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries unmanaged address (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:154 assert (address_ok, \"'B' channel PutFull carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries source that is not first source (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:155 assert (legal_source, \"'B' channel PutFull carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:156 assert (is_aligned, \"'B' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries invalid param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:157 assert (bundle.param === UInt(0), \"'B' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull contains invalid mask (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:158 assert (bundle.mask === mask, \"'B' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutPartial type unsupported by client (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:162 assert (edge.client.supportsPutPartial(bundle.source, bundle.size), \"'B' channel carries PutPartial type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:163 assert (address_ok, \"'B' channel PutPartial carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:164 assert (legal_source, \"'B' channel PutPartial carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:165 assert (is_aligned, \"'B' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries invalid param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:166 assert (bundle.param === UInt(0), \"'B' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial contains invalid mask (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:167 assert ((bundle.mask & ~mask) === UInt(0), \"'B' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Arithmetic type unsupported by client (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:171 assert (edge.client.supportsArithmetic(bundle.source, bundle.size), \"'B' channel carries Arithmetic type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:172 assert (address_ok, \"'B' channel Arithmetic carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:173 assert (legal_source, \"'B' channel Arithmetic carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:174 assert (is_aligned, \"'B' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries invalid opcode param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:175 assert (TLAtomics.isArithmetic(bundle.param), \"'B' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:176 assert (bundle.mask === mask, \"'B' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Logical type unsupported by client (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:180 assert (edge.client.supportsLogical(bundle.source, bundle.size), \"'B' channel carries Logical type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries unmanaged address (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:181 assert (address_ok, \"'B' channel Logical carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries source that is not first source (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:182 assert (legal_source, \"'B' channel Logical carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:183 assert (is_aligned, \"'B' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries invalid opcode param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:184 assert (TLAtomics.isLogical(bundle.param), \"'B' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical contains invalid mask (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:185 assert (bundle.mask === mask, \"'B' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Hint type unsupported by client (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:189 assert (edge.client.supportsHint(bundle.source, bundle.size), \"'B' channel carries Hint type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries unmanaged address (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:190 assert (address_ok, \"'B' channel Hint carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries source that is not first source (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:191 assert (legal_source, \"'B' channel Hint carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:192 assert (is_aligned, \"'B' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint contains invalid mask (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:193 assert (bundle.mask === mask, \"'B' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint is corrupt (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:194 assert (!bundle.corrupt, \"'B' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel has invalid opcode (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:199 assert (TLMessages.isC(bundle.opcode), \"'C' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:205 assert (visible(edge.address(bundle), bundle.source, edge), \"'C' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1807) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:208 assert (address_ok, \"'C' channel ProbeAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1807) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1810) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:209 assert (source_ok, \"'C' channel ProbeAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1810) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1814) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:210 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1814) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1817) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:211 assert (is_aligned, \"'C' channel ProbeAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1817) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1821) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:212 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAck carries invalid report param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1821) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1825) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck is corrupt (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:213 assert (!bundle.corrupt, \"'C' channel ProbeAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1825) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_187 & _T_1807) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:217 assert (address_ok, \"'C' channel ProbeAckData carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_187 & _T_1807) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_187 & _T_1810) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:218 assert (source_ok, \"'C' channel ProbeAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_187 & _T_1810) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_187 & _T_1814) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:219 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAckData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_187 & _T_1814) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_187 & _T_1817) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:220 assert (is_aligned, \"'C' channel ProbeAckData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_187 & _T_1817) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_187 & _T_1821) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:221 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAckData carries invalid report param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_187 & _T_1821) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1872) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:225 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries Release type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1872) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1959) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:226 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1959) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1810) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:227 assert (source_ok, \"'C' channel Release carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1810) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1814) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:228 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel Release smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1814) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1817) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:229 assert (is_aligned, \"'C' channel Release address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1817) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1973) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid shrink param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:230 assert (TLPermissions.isShrink(bundle.param), \"'C' channel Release carries invalid shrink param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1973) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1825) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release is corrupt (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:231 assert (!bundle.corrupt, \"'C' channel Release is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1825) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1872) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:235 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries ReleaseData type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1872) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1959) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:236 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1959) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1810) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:237 assert (source_ok, \"'C' channel ReleaseData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1810) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1814) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:238 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ReleaseData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1814) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1817) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:239 assert (is_aligned, \"'C' channel ReleaseData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1817) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1973) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid shrink param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:240 assert (TLPermissions.isShrink(bundle.param), \"'C' channel ReleaseData carries invalid shrink param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1973) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_1807) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:244 assert (address_ok, \"'C' channel AccessAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_1807) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_1810) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:245 assert (source_ok, \"'C' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_1810) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_1817) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:246 assert (is_aligned, \"'C' channel AccessAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_1817) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_2121) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:247 assert (bundle.param === UInt(0), \"'C' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_2121) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_1825) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck is corrupt (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:248 assert (!bundle.corrupt, \"'C' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_1825) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_1807) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:252 assert (address_ok, \"'C' channel AccessAckData carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_1807) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_1810) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:253 assert (source_ok, \"'C' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_1810) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_1817) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:254 assert (is_aligned, \"'C' channel AccessAckData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_1817) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_2121) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:255 assert (bundle.param === UInt(0), \"'C' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_2121) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1807) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:259 assert (address_ok, \"'C' channel HintAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1807) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1810) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:260 assert (source_ok, \"'C' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1810) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1817) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:261 assert (is_aligned, \"'C' channel HintAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1817) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_2121) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:262 assert (bundle.param === UInt(0), \"'C' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_2121) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1825) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck is corrupt (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:263 assert (!bundle.corrupt, \"'C' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1825) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_e_valid & _T_2161) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channels carries invalid sink ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:330 assert (sink_ok, \"'E' channels carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_e_valid & _T_2161) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2188 & _T_2192) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2188 & _T_2192) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2188 & _T_2196) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2188 & _T_2196) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2188 & _T_2200) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2188 & _T_2200) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2188 & _T_2204) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2188 & _T_2204) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2188 & _T_2208) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2188 & _T_2208) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2237 & _T_2241) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2237 & _T_2241) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2237 & _T_2245) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2237 & _T_2245) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2237 & _T_2249) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2237 & _T_2249) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2237 & _T_2253) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2237 & _T_2253) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2237 & _T_2257) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2237 & _T_2257) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2237 & _T_2261) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2237 & _T_2261) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:378 assert (b.bits.opcode === opcode, \"'B' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:379 assert (b.bits.param  === param,  \"'B' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel size changed within multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:380 assert (b.bits.size   === size,   \"'B' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel source changed within multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:381 assert (b.bits.source === source, \"'B' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:382 assert (b.bits.address=== address,\"'B' channel addresss changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2338 & _T_2342) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:401 assert (c.bits.opcode === opcode, \"'C' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2338 & _T_2342) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2338 & _T_2346) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:402 assert (c.bits.param  === param,  \"'C' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2338 & _T_2346) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2338 & _T_2350) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:403 assert (c.bits.size   === size,   \"'C' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2338 & _T_2350) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2338 & _T_2354) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:404 assert (c.bits.source === source, \"'C' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2338 & _T_2354) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2338 & _T_2358) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:405 assert (c.bits.address=== address,\"'C' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2338 & _T_2358) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2403 & _T_2411) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2403 & _T_2411) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2418 & _T_2425) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2418 & _T_2425) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2432) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2432) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2445) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:479 assert (!inflight.orR || limit === UInt(0) || watchdog < limit, \"TileLink timeout expired\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2445) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2478 & _T_2485) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:494 assert(!inflight(bundle.d.bits.sink), \"'D' channel re-used a sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2478 & _T_2485) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2487 & _T_2496) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at ChiplinkTest.scala:362:47)\n    at Monitor.scala:500 assert((d_set | inflight)(bundle.e.bits.sink), \"'E' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2487 & _T_2496) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLMonitor_15( 
  input         clock, 
  input         reset, 
  input         io_in_a_ready, 
  input         io_in_a_valid, 
  input  [2:0]  io_in_a_bits_opcode, 
  input  [2:0]  io_in_a_bits_param, 
  input  [3:0]  io_in_a_bits_size, 
  input  [6:0]  io_in_a_bits_source, 
  input  [31:0] io_in_a_bits_address, 
  input  [7:0]  io_in_a_bits_mask, 
  input         io_in_c_ready, 
  input         io_in_c_valid, 
  input  [2:0]  io_in_c_bits_opcode, 
  input  [2:0]  io_in_c_bits_param, 
  input  [3:0]  io_in_c_bits_size, 
  input  [6:0]  io_in_c_bits_source, 
  input  [31:0] io_in_c_bits_address, 
  input         io_in_c_bits_corrupt, 
  input         io_in_d_ready, 
  input         io_in_d_valid, 
  input  [2:0]  io_in_d_bits_opcode, 
  input  [1:0]  io_in_d_bits_param, 
  input  [3:0]  io_in_d_bits_size, 
  input  [6:0]  io_in_d_bits_source, 
  input         io_in_d_bits_sink, 
  input         io_in_d_bits_denied, 
  input         io_in_d_bits_corrupt, 
  input         io_in_e_ready, 
  input         io_in_e_valid, 
  input         io_in_e_bits_sink 
);
  wire [31:0] plusarg_reader_out; 
  wire [2:0] _T_7; 
  wire  _T_8; 
  wire  _T_16; 
  wire  _T_24; 
  wire  _T_32; 
  wire  _T_40; 
  wire  _T_48; 
  wire  _T_56; 
  wire  _T_64; 
  wire  _T_70; 
  wire  _T_71; 
  wire  _T_72; 
  wire  _T_73; 
  wire  _T_74; 
  wire  _T_75; 
  wire  _T_76; 
  wire [22:0] _T_78; 
  wire [7:0] _T_79; 
  wire [7:0] _T_80; 
  wire [31:0] _GEN_33; 
  wire [31:0] _T_81; 
  wire  _T_82; 
  wire [1:0] _T_84; 
  wire [3:0] _T_85; 
  wire [2:0] _T_86; 
  wire [2:0] _T_87; 
  wire  _T_88; 
  wire  _T_89; 
  wire  _T_90; 
  wire  _T_91; 
  wire  _T_93; 
  wire  _T_94; 
  wire  _T_96; 
  wire  _T_97; 
  wire  _T_98; 
  wire  _T_99; 
  wire  _T_100; 
  wire  _T_101; 
  wire  _T_102; 
  wire  _T_103; 
  wire  _T_104; 
  wire  _T_105; 
  wire  _T_106; 
  wire  _T_107; 
  wire  _T_108; 
  wire  _T_109; 
  wire  _T_110; 
  wire  _T_111; 
  wire  _T_112; 
  wire  _T_113; 
  wire  _T_114; 
  wire  _T_115; 
  wire  _T_116; 
  wire  _T_117; 
  wire  _T_118; 
  wire  _T_119; 
  wire  _T_120; 
  wire  _T_121; 
  wire  _T_122; 
  wire  _T_123; 
  wire  _T_124; 
  wire  _T_125; 
  wire  _T_126; 
  wire  _T_127; 
  wire  _T_128; 
  wire  _T_129; 
  wire  _T_130; 
  wire  _T_131; 
  wire  _T_132; 
  wire  _T_133; 
  wire  _T_134; 
  wire  _T_135; 
  wire  _T_136; 
  wire  _T_137; 
  wire  _T_138; 
  wire  _T_139; 
  wire [7:0] _T_146; 
  wire  _T_277; 
  wire [31:0] _T_279; 
  wire [32:0] _T_280; 
  wire [32:0] _T_281; 
  wire [32:0] _T_282; 
  wire  _T_283; 
  wire [31:0] _T_284; 
  wire [32:0] _T_285; 
  wire [32:0] _T_286; 
  wire [32:0] _T_287; 
  wire  _T_288; 
  wire  _T_289; 
  wire  _T_292; 
  wire [31:0] _T_295; 
  wire [32:0] _T_296; 
  wire [32:0] _T_297; 
  wire [32:0] _T_298; 
  wire  _T_299; 
  wire  _T_300; 
  wire  _T_304; 
  wire  _T_305; 
  wire  _T_374; 
  wire  _T_391; 
  wire  _T_392; 
  wire  _T_394; 
  wire  _T_395; 
  wire  _T_398; 
  wire  _T_399; 
  wire  _T_401; 
  wire  _T_402; 
  wire  _T_403; 
  wire  _T_405; 
  wire  _T_406; 
  wire [7:0] _T_407; 
  wire  _T_408; 
  wire  _T_410; 
  wire  _T_411; 
  wire  _T_416; 
  wire  _T_546; 
  wire  _T_548; 
  wire  _T_549; 
  wire  _T_559; 
  wire  _T_580; 
  wire  _T_581; 
  wire  _T_584; 
  wire  _T_585; 
  wire  _T_592; 
  wire  _T_594; 
  wire  _T_595; 
  wire  _T_596; 
  wire  _T_598; 
  wire  _T_599; 
  wire  _T_604; 
  wire  _T_619; 
  wire  _T_620; 
  wire  _T_622; 
  wire  _T_630; 
  wire  _T_632; 
  wire  _T_634; 
  wire  _T_635; 
  wire  _T_650; 
  wire [7:0] _T_692; 
  wire [7:0] _T_693; 
  wire  _T_694; 
  wire  _T_696; 
  wire  _T_697; 
  wire  _T_698; 
  wire  _T_700; 
  wire  _T_720; 
  wire  _T_723; 
  wire  _T_724; 
  wire  _T_731; 
  wire  _T_733; 
  wire  _T_734; 
  wire  _T_739; 
  wire  _T_772; 
  wire  _T_774; 
  wire  _T_775; 
  wire  _T_780; 
  wire  _T_823; 
  wire  _T_825; 
  wire  _T_826; 
  wire [2:0] _T_829; 
  wire  _T_830; 
  wire  _T_838; 
  wire  _T_846; 
  wire  _T_854; 
  wire  _T_862; 
  wire  _T_870; 
  wire  _T_878; 
  wire  _T_886; 
  wire  _T_892; 
  wire  _T_893; 
  wire  _T_894; 
  wire  _T_895; 
  wire  _T_896; 
  wire  _T_897; 
  wire  _T_898; 
  wire  _T_899; 
  wire  _T_900; 
  wire  _T_902; 
  wire  _T_903; 
  wire  _T_904; 
  wire  _T_906; 
  wire  _T_907; 
  wire  _T_908; 
  wire  _T_910; 
  wire  _T_911; 
  wire  _T_912; 
  wire  _T_914; 
  wire  _T_915; 
  wire  _T_916; 
  wire  _T_918; 
  wire  _T_919; 
  wire  _T_920; 
  wire  _T_925; 
  wire  _T_926; 
  wire  _T_931; 
  wire  _T_933; 
  wire  _T_934; 
  wire  _T_935; 
  wire  _T_937; 
  wire  _T_938; 
  wire  _T_948; 
  wire  _T_968; 
  wire  _T_970; 
  wire  _T_971; 
  wire  _T_977; 
  wire  _T_994; 
  wire  _T_1012; 
  wire [2:0] _T_1580; 
  wire  _T_1581; 
  wire  _T_1589; 
  wire  _T_1597; 
  wire  _T_1605; 
  wire  _T_1613; 
  wire  _T_1621; 
  wire  _T_1629; 
  wire  _T_1637; 
  wire  _T_1643; 
  wire  _T_1644; 
  wire  _T_1645; 
  wire  _T_1646; 
  wire  _T_1647; 
  wire  _T_1648; 
  wire  _T_1649; 
  wire [22:0] _T_1651; 
  wire [7:0] _T_1652; 
  wire [7:0] _T_1653; 
  wire [31:0] _GEN_34; 
  wire [31:0] _T_1654; 
  wire  _T_1655; 
  wire [31:0] _T_1656; 
  wire [32:0] _T_1657; 
  wire [32:0] _T_1658; 
  wire [32:0] _T_1659; 
  wire  _T_1660; 
  wire [31:0] _T_1661; 
  wire [32:0] _T_1662; 
  wire [32:0] _T_1663; 
  wire [32:0] _T_1664; 
  wire  _T_1665; 
  wire [31:0] _T_1666; 
  wire [32:0] _T_1667; 
  wire [32:0] _T_1668; 
  wire [32:0] _T_1669; 
  wire  _T_1670; 
  wire  _T_1672; 
  wire  _T_1673; 
  wire  _T_1804; 
  wire  _T_1806; 
  wire  _T_1807; 
  wire  _T_1809; 
  wire  _T_1810; 
  wire  _T_1811; 
  wire  _T_1813; 
  wire  _T_1814; 
  wire  _T_1816; 
  wire  _T_1817; 
  wire  _T_1818; 
  wire  _T_1820; 
  wire  _T_1821; 
  wire  _T_1822; 
  wire  _T_1824; 
  wire  _T_1825; 
  wire  _T_1826; 
  wire  _T_1844; 
  wire  _T_1859; 
  wire  _T_1867; 
  wire  _T_1871; 
  wire  _T_1872; 
  wire  _T_1941; 
  wire  _T_1958; 
  wire  _T_1959; 
  wire  _T_1970; 
  wire  _T_1972; 
  wire  _T_1973; 
  wire  _T_1978; 
  wire  _T_2108; 
  wire  _T_2118; 
  wire  _T_2120; 
  wire  _T_2121; 
  wire  _T_2126; 
  wire  _T_2140; 
  wire  _T_2158; 
  wire  _T_2160; 
  wire  _T_2161; 
  wire  _T_2162; 
  wire [4:0] _T_2167; 
  wire  _T_2168; 
  wire  _T_2169; 
  reg [4:0] _T_2171; 
  reg [31:0] _RAND_0;
  wire [4:0] _T_2173; 
  wire  _T_2174; 
  reg [2:0] _T_2182; 
  reg [31:0] _RAND_1;
  reg [2:0] _T_2183; 
  reg [31:0] _RAND_2;
  reg [3:0] _T_2184; 
  reg [31:0] _RAND_3;
  reg [6:0] _T_2185; 
  reg [31:0] _RAND_4;
  reg [31:0] _T_2186; 
  reg [31:0] _RAND_5;
  wire  _T_2187; 
  wire  _T_2188; 
  wire  _T_2189; 
  wire  _T_2191; 
  wire  _T_2192; 
  wire  _T_2193; 
  wire  _T_2195; 
  wire  _T_2196; 
  wire  _T_2197; 
  wire  _T_2199; 
  wire  _T_2200; 
  wire  _T_2201; 
  wire  _T_2203; 
  wire  _T_2204; 
  wire  _T_2205; 
  wire  _T_2207; 
  wire  _T_2208; 
  wire  _T_2210; 
  wire  _T_2211; 
  wire [22:0] _T_2213; 
  wire [7:0] _T_2214; 
  wire [7:0] _T_2215; 
  wire [4:0] _T_2216; 
  wire  _T_2217; 
  reg [4:0] _T_2219; 
  reg [31:0] _RAND_6;
  wire [4:0] _T_2221; 
  wire  _T_2222; 
  reg [2:0] _T_2230; 
  reg [31:0] _RAND_7;
  reg [1:0] _T_2231; 
  reg [31:0] _RAND_8;
  reg [3:0] _T_2232; 
  reg [31:0] _RAND_9;
  reg [6:0] _T_2233; 
  reg [31:0] _RAND_10;
  reg  _T_2234; 
  reg [31:0] _RAND_11;
  reg  _T_2235; 
  reg [31:0] _RAND_12;
  wire  _T_2236; 
  wire  _T_2237; 
  wire  _T_2238; 
  wire  _T_2240; 
  wire  _T_2241; 
  wire  _T_2242; 
  wire  _T_2244; 
  wire  _T_2245; 
  wire  _T_2246; 
  wire  _T_2248; 
  wire  _T_2249; 
  wire  _T_2250; 
  wire  _T_2252; 
  wire  _T_2253; 
  wire  _T_2254; 
  wire  _T_2256; 
  wire  _T_2257; 
  wire  _T_2258; 
  wire  _T_2260; 
  wire  _T_2261; 
  wire  _T_2263; 
  wire  _T_2313; 
  wire [4:0] _T_2318; 
  wire  _T_2319; 
  reg [4:0] _T_2321; 
  reg [31:0] _RAND_13;
  wire [4:0] _T_2323; 
  wire  _T_2324; 
  reg [2:0] _T_2332; 
  reg [31:0] _RAND_14;
  reg [2:0] _T_2333; 
  reg [31:0] _RAND_15;
  reg [3:0] _T_2334; 
  reg [31:0] _RAND_16;
  reg [6:0] _T_2335; 
  reg [31:0] _RAND_17;
  reg [31:0] _T_2336; 
  reg [31:0] _RAND_18;
  wire  _T_2337; 
  wire  _T_2338; 
  wire  _T_2339; 
  wire  _T_2341; 
  wire  _T_2342; 
  wire  _T_2343; 
  wire  _T_2345; 
  wire  _T_2346; 
  wire  _T_2347; 
  wire  _T_2349; 
  wire  _T_2350; 
  wire  _T_2351; 
  wire  _T_2353; 
  wire  _T_2354; 
  wire  _T_2355; 
  wire  _T_2357; 
  wire  _T_2358; 
  wire  _T_2360; 
  reg [127:0] _T_2361; 
  reg [127:0] _RAND_19;
  reg [4:0] _T_2371; 
  reg [31:0] _RAND_20;
  wire [4:0] _T_2373; 
  wire  _T_2374; 
  reg [4:0] _T_2390; 
  reg [31:0] _RAND_21;
  wire [4:0] _T_2392; 
  wire  _T_2393; 
  wire  _T_2403; 
  wire [127:0] _T_2405; 
  wire [127:0] _T_2406; 
  wire  _T_2407; 
  wire  _T_2408; 
  wire  _T_2410; 
  wire  _T_2411; 
  wire [127:0] _GEN_27; 
  wire  _T_2415; 
  wire  _T_2417; 
  wire  _T_2418; 
  wire [127:0] _T_2419; 
  wire [127:0] _T_2420; 
  wire [127:0] _T_2421; 
  wire  _T_2422; 
  wire  _T_2424; 
  wire  _T_2425; 
  wire [127:0] _GEN_28; 
  wire  _T_2426; 
  wire  _T_2427; 
  wire  _T_2428; 
  wire  _T_2429; 
  wire  _T_2431; 
  wire  _T_2432; 
  wire [127:0] _T_2433; 
  wire [127:0] _T_2434; 
  wire [127:0] _T_2435; 
  reg [31:0] _T_2436; 
  reg [31:0] _RAND_22;
  wire  _T_2437; 
  wire  _T_2438; 
  wire  _T_2439; 
  wire  _T_2440; 
  wire  _T_2441; 
  wire  _T_2442; 
  wire  _T_2444; 
  wire  _T_2445; 
  wire [31:0] _T_2447; 
  wire  _T_2450; 
  reg  _T_2451; 
  reg [31:0] _RAND_23;
  reg [4:0] _T_2460; 
  reg [31:0] _RAND_24;
  wire [4:0] _T_2462; 
  wire  _T_2463; 
  wire  _T_2473; 
  wire  _T_2474; 
  wire  _T_2475; 
  wire  _T_2476; 
  wire  _T_2477; 
  wire  _T_2478; 
  wire [1:0] _T_2479; 
  wire  _T_2480; 
  wire  _T_2482; 
  wire  _T_2484; 
  wire  _T_2485; 
  wire [1:0] _GEN_31; 
  wire  _T_2487; 
  wire [1:0] _T_2490; 
  wire  _T_2471; 
  wire  _T_2491; 
  wire  _T_2492; 
  wire  _T_2495; 
  wire  _T_2496; 
  wire [1:0] _GEN_32; 
  wire  _T_2497; 
  wire  _T_2486; 
  wire  _T_2498; 
  wire  _T_2499; 
  wire  _GEN_35; 
  wire  _GEN_49; 
  wire  _GEN_65; 
  wire  _GEN_75; 
  wire  _GEN_85; 
  wire  _GEN_95; 
  wire  _GEN_105; 
  wire  _GEN_115; 
  wire  _GEN_123; 
  wire  _GEN_133; 
  wire  _GEN_145; 
  wire  _GEN_157; 
  wire  _GEN_163; 
  wire  _GEN_169; 
  wire  _GEN_175; 
  wire  _GEN_187; 
  wire  _GEN_197; 
  wire  _GEN_211; 
  wire  _GEN_223; 
  wire  _GEN_233; 
  wire  _GEN_241; 
  dual_plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0)) plusarg_reader ( 
    .out(plusarg_reader_out)
  );
  assign _T_7 = io_in_a_bits_source[6:4]; 
  assign _T_8 = _T_7 == 3'h0; 
  assign _T_16 = _T_7 == 3'h1; 
  assign _T_24 = _T_7 == 3'h2; 
  assign _T_32 = _T_7 == 3'h3; 
  assign _T_40 = _T_7 == 3'h4; 
  assign _T_48 = _T_7 == 3'h5; 
  assign _T_56 = _T_7 == 3'h6; 
  assign _T_64 = _T_7 == 3'h7; 
  assign _T_70 = _T_8 | _T_16; 
  assign _T_71 = _T_70 | _T_24; 
  assign _T_72 = _T_71 | _T_32; 
  assign _T_73 = _T_72 | _T_40; 
  assign _T_74 = _T_73 | _T_48; 
  assign _T_75 = _T_74 | _T_56; 
  assign _T_76 = _T_75 | _T_64; 
  assign _T_78 = 23'hff << io_in_a_bits_size; 
  assign _T_79 = _T_78[7:0]; 
  assign _T_80 = ~ _T_79; 
  assign _GEN_33 = {{24'd0}, _T_80}; 
  assign _T_81 = io_in_a_bits_address & _GEN_33; 
  assign _T_82 = _T_81 == 32'h0; 
  assign _T_84 = io_in_a_bits_size[1:0]; 
  assign _T_85 = 4'h1 << _T_84; 
  assign _T_86 = _T_85[2:0]; 
  assign _T_87 = _T_86 | 3'h1; 
  assign _T_88 = io_in_a_bits_size >= 4'h3; 
  assign _T_89 = _T_87[2]; 
  assign _T_90 = io_in_a_bits_address[2]; 
  assign _T_91 = _T_90 == 1'h0; 
  assign _T_93 = _T_89 & _T_91; 
  assign _T_94 = _T_88 | _T_93; 
  assign _T_96 = _T_89 & _T_90; 
  assign _T_97 = _T_88 | _T_96; 
  assign _T_98 = _T_87[1]; 
  assign _T_99 = io_in_a_bits_address[1]; 
  assign _T_100 = _T_99 == 1'h0; 
  assign _T_101 = _T_91 & _T_100; 
  assign _T_102 = _T_98 & _T_101; 
  assign _T_103 = _T_94 | _T_102; 
  assign _T_104 = _T_91 & _T_99; 
  assign _T_105 = _T_98 & _T_104; 
  assign _T_106 = _T_94 | _T_105; 
  assign _T_107 = _T_90 & _T_100; 
  assign _T_108 = _T_98 & _T_107; 
  assign _T_109 = _T_97 | _T_108; 
  assign _T_110 = _T_90 & _T_99; 
  assign _T_111 = _T_98 & _T_110; 
  assign _T_112 = _T_97 | _T_111; 
  assign _T_113 = _T_87[0]; 
  assign _T_114 = io_in_a_bits_address[0]; 
  assign _T_115 = _T_114 == 1'h0; 
  assign _T_116 = _T_101 & _T_115; 
  assign _T_117 = _T_113 & _T_116; 
  assign _T_118 = _T_103 | _T_117; 
  assign _T_119 = _T_101 & _T_114; 
  assign _T_120 = _T_113 & _T_119; 
  assign _T_121 = _T_103 | _T_120; 
  assign _T_122 = _T_104 & _T_115; 
  assign _T_123 = _T_113 & _T_122; 
  assign _T_124 = _T_106 | _T_123; 
  assign _T_125 = _T_104 & _T_114; 
  assign _T_126 = _T_113 & _T_125; 
  assign _T_127 = _T_106 | _T_126; 
  assign _T_128 = _T_107 & _T_115; 
  assign _T_129 = _T_113 & _T_128; 
  assign _T_130 = _T_109 | _T_129; 
  assign _T_131 = _T_107 & _T_114; 
  assign _T_132 = _T_113 & _T_131; 
  assign _T_133 = _T_109 | _T_132; 
  assign _T_134 = _T_110 & _T_115; 
  assign _T_135 = _T_113 & _T_134; 
  assign _T_136 = _T_112 | _T_135; 
  assign _T_137 = _T_110 & _T_114; 
  assign _T_138 = _T_113 & _T_137; 
  assign _T_139 = _T_112 | _T_138; 
  assign _T_146 = {_T_139,_T_136,_T_133,_T_130,_T_127,_T_124,_T_121,_T_118}; 
  assign _T_277 = io_in_a_bits_opcode == 3'h6; 
  assign _T_279 = io_in_a_bits_address ^ 32'h80000000; 
  assign _T_280 = {1'b0,$signed(_T_279)}; 
  assign _T_281 = $signed(_T_280) & $signed(-33'sh80000000); 
  assign _T_282 = $signed(_T_281); 
  assign _T_283 = $signed(_T_282) == $signed(33'sh0); 
  assign _T_284 = io_in_a_bits_address ^ 32'h40000000; 
  assign _T_285 = {1'b0,$signed(_T_284)}; 
  assign _T_286 = $signed(_T_285) & $signed(-33'sh20000000); 
  assign _T_287 = $signed(_T_286); 
  assign _T_288 = $signed(_T_287) == $signed(33'sh0); 
  assign _T_289 = _T_283 | _T_288; 
  assign _T_292 = io_in_a_bits_size <= 4'h6; 
  assign _T_295 = io_in_a_bits_address ^ 32'h10000000; 
  assign _T_296 = {1'b0,$signed(_T_295)}; 
  assign _T_297 = $signed(_T_296) & $signed(-33'sh10000000); 
  assign _T_298 = $signed(_T_297); 
  assign _T_299 = $signed(_T_298) == $signed(33'sh0); 
  assign _T_300 = _T_292 & _T_299; 
  assign _T_304 = _T_300 | reset; 
  assign _T_305 = _T_304 == 1'h0; 
  assign _T_374 = _T_8 ? _T_292 : 1'h0; 
  assign _T_391 = _T_374 | reset; 
  assign _T_392 = _T_391 == 1'h0; 
  assign _T_394 = _T_76 | reset; 
  assign _T_395 = _T_394 == 1'h0; 
  assign _T_398 = _T_88 | reset; 
  assign _T_399 = _T_398 == 1'h0; 
  assign _T_401 = _T_82 | reset; 
  assign _T_402 = _T_401 == 1'h0; 
  assign _T_403 = io_in_a_bits_param <= 3'h2; 
  assign _T_405 = _T_403 | reset; 
  assign _T_406 = _T_405 == 1'h0; 
  assign _T_407 = ~ io_in_a_bits_mask; 
  assign _T_408 = _T_407 == 8'h0; 
  assign _T_410 = _T_408 | reset; 
  assign _T_411 = _T_410 == 1'h0; 
  assign _T_416 = io_in_a_bits_opcode == 3'h7; 
  assign _T_546 = io_in_a_bits_param != 3'h0; 
  assign _T_548 = _T_546 | reset; 
  assign _T_549 = _T_548 == 1'h0; 
  assign _T_559 = io_in_a_bits_opcode == 3'h4; 
  assign _T_580 = _T_289 | _T_299; 
  assign _T_581 = _T_292 & _T_580; 
  assign _T_584 = _T_581 | reset; 
  assign _T_585 = _T_584 == 1'h0; 
  assign _T_592 = io_in_a_bits_param == 3'h0; 
  assign _T_594 = _T_592 | reset; 
  assign _T_595 = _T_594 == 1'h0; 
  assign _T_596 = io_in_a_bits_mask == _T_146; 
  assign _T_598 = _T_596 | reset; 
  assign _T_599 = _T_598 == 1'h0; 
  assign _T_604 = io_in_a_bits_opcode == 3'h0; 
  assign _T_619 = _T_283 | _T_299; 
  assign _T_620 = _T_292 & _T_619; 
  assign _T_622 = io_in_a_bits_size <= 4'h8; 
  assign _T_630 = _T_622 & _T_288; 
  assign _T_632 = _T_620 | _T_630; 
  assign _T_634 = _T_632 | reset; 
  assign _T_635 = _T_634 == 1'h0; 
  assign _T_650 = io_in_a_bits_opcode == 3'h1; 
  assign _T_692 = ~ _T_146; 
  assign _T_693 = io_in_a_bits_mask & _T_692; 
  assign _T_694 = _T_693 == 8'h0; 
  assign _T_696 = _T_694 | reset; 
  assign _T_697 = _T_696 == 1'h0; 
  assign _T_698 = io_in_a_bits_opcode == 3'h2; 
  assign _T_700 = io_in_a_bits_size <= 4'h3; 
  assign _T_720 = _T_700 & _T_580; 
  assign _T_723 = _T_720 | reset; 
  assign _T_724 = _T_723 == 1'h0; 
  assign _T_731 = io_in_a_bits_param <= 3'h4; 
  assign _T_733 = _T_731 | reset; 
  assign _T_734 = _T_733 == 1'h0; 
  assign _T_739 = io_in_a_bits_opcode == 3'h3; 
  assign _T_772 = io_in_a_bits_param <= 3'h3; 
  assign _T_774 = _T_772 | reset; 
  assign _T_775 = _T_774 == 1'h0; 
  assign _T_780 = io_in_a_bits_opcode == 3'h5; 
  assign _T_823 = io_in_d_bits_opcode <= 3'h6; 
  assign _T_825 = _T_823 | reset; 
  assign _T_826 = _T_825 == 1'h0; 
  assign _T_829 = io_in_d_bits_source[6:4]; 
  assign _T_830 = _T_829 == 3'h0; 
  assign _T_838 = _T_829 == 3'h1; 
  assign _T_846 = _T_829 == 3'h2; 
  assign _T_854 = _T_829 == 3'h3; 
  assign _T_862 = _T_829 == 3'h4; 
  assign _T_870 = _T_829 == 3'h5; 
  assign _T_878 = _T_829 == 3'h6; 
  assign _T_886 = _T_829 == 3'h7; 
  assign _T_892 = _T_830 | _T_838; 
  assign _T_893 = _T_892 | _T_846; 
  assign _T_894 = _T_893 | _T_854; 
  assign _T_895 = _T_894 | _T_862; 
  assign _T_896 = _T_895 | _T_870; 
  assign _T_897 = _T_896 | _T_878; 
  assign _T_898 = _T_897 | _T_886; 
  assign _T_899 = io_in_d_bits_sink < 1'h1; 
  assign _T_900 = io_in_d_bits_opcode == 3'h6; 
  assign _T_902 = _T_898 | reset; 
  assign _T_903 = _T_902 == 1'h0; 
  assign _T_904 = io_in_d_bits_size >= 4'h3; 
  assign _T_906 = _T_904 | reset; 
  assign _T_907 = _T_906 == 1'h0; 
  assign _T_908 = io_in_d_bits_param == 2'h0; 
  assign _T_910 = _T_908 | reset; 
  assign _T_911 = _T_910 == 1'h0; 
  assign _T_912 = io_in_d_bits_corrupt == 1'h0; 
  assign _T_914 = _T_912 | reset; 
  assign _T_915 = _T_914 == 1'h0; 
  assign _T_916 = io_in_d_bits_denied == 1'h0; 
  assign _T_918 = _T_916 | reset; 
  assign _T_919 = _T_918 == 1'h0; 
  assign _T_920 = io_in_d_bits_opcode == 3'h4; 
  assign _T_925 = _T_899 | reset; 
  assign _T_926 = _T_925 == 1'h0; 
  assign _T_931 = io_in_d_bits_param <= 2'h2; 
  assign _T_933 = _T_931 | reset; 
  assign _T_934 = _T_933 == 1'h0; 
  assign _T_935 = io_in_d_bits_param != 2'h2; 
  assign _T_937 = _T_935 | reset; 
  assign _T_938 = _T_937 == 1'h0; 
  assign _T_948 = io_in_d_bits_opcode == 3'h5; 
  assign _T_968 = _T_916 | io_in_d_bits_corrupt; 
  assign _T_970 = _T_968 | reset; 
  assign _T_971 = _T_970 == 1'h0; 
  assign _T_977 = io_in_d_bits_opcode == 3'h0; 
  assign _T_994 = io_in_d_bits_opcode == 3'h1; 
  assign _T_1012 = io_in_d_bits_opcode == 3'h2; 
  assign _T_1580 = io_in_c_bits_source[6:4]; 
  assign _T_1581 = _T_1580 == 3'h0; 
  assign _T_1589 = _T_1580 == 3'h1; 
  assign _T_1597 = _T_1580 == 3'h2; 
  assign _T_1605 = _T_1580 == 3'h3; 
  assign _T_1613 = _T_1580 == 3'h4; 
  assign _T_1621 = _T_1580 == 3'h5; 
  assign _T_1629 = _T_1580 == 3'h6; 
  assign _T_1637 = _T_1580 == 3'h7; 
  assign _T_1643 = _T_1581 | _T_1589; 
  assign _T_1644 = _T_1643 | _T_1597; 
  assign _T_1645 = _T_1644 | _T_1605; 
  assign _T_1646 = _T_1645 | _T_1613; 
  assign _T_1647 = _T_1646 | _T_1621; 
  assign _T_1648 = _T_1647 | _T_1629; 
  assign _T_1649 = _T_1648 | _T_1637; 
  assign _T_1651 = 23'hff << io_in_c_bits_size; 
  assign _T_1652 = _T_1651[7:0]; 
  assign _T_1653 = ~ _T_1652; 
  assign _GEN_34 = {{24'd0}, _T_1653}; 
  assign _T_1654 = io_in_c_bits_address & _GEN_34; 
  assign _T_1655 = _T_1654 == 32'h0; 
  assign _T_1656 = io_in_c_bits_address ^ 32'h80000000; 
  assign _T_1657 = {1'b0,$signed(_T_1656)}; 
  assign _T_1658 = $signed(_T_1657) & $signed(-33'sh80000000); 
  assign _T_1659 = $signed(_T_1658); 
  assign _T_1660 = $signed(_T_1659) == $signed(33'sh0); 
  assign _T_1661 = io_in_c_bits_address ^ 32'h40000000; 
  assign _T_1662 = {1'b0,$signed(_T_1661)}; 
  assign _T_1663 = $signed(_T_1662) & $signed(-33'sh20000000); 
  assign _T_1664 = $signed(_T_1663); 
  assign _T_1665 = $signed(_T_1664) == $signed(33'sh0); 
  assign _T_1666 = io_in_c_bits_address ^ 32'h10000000; 
  assign _T_1667 = {1'b0,$signed(_T_1666)}; 
  assign _T_1668 = $signed(_T_1667) & $signed(-33'sh10000000); 
  assign _T_1669 = $signed(_T_1668); 
  assign _T_1670 = $signed(_T_1669) == $signed(33'sh0); 
  assign _T_1672 = _T_1660 | _T_1665; 
  assign _T_1673 = _T_1672 | _T_1670; 
  assign _T_1804 = io_in_c_bits_opcode == 3'h4; 
  assign _T_1806 = _T_1673 | reset; 
  assign _T_1807 = _T_1806 == 1'h0; 
  assign _T_1809 = _T_1649 | reset; 
  assign _T_1810 = _T_1809 == 1'h0; 
  assign _T_1811 = io_in_c_bits_size >= 4'h3; 
  assign _T_1813 = _T_1811 | reset; 
  assign _T_1814 = _T_1813 == 1'h0; 
  assign _T_1816 = _T_1655 | reset; 
  assign _T_1817 = _T_1816 == 1'h0; 
  assign _T_1818 = io_in_c_bits_param <= 3'h5; 
  assign _T_1820 = _T_1818 | reset; 
  assign _T_1821 = _T_1820 == 1'h0; 
  assign _T_1822 = io_in_c_bits_corrupt == 1'h0; 
  assign _T_1824 = _T_1822 | reset; 
  assign _T_1825 = _T_1824 == 1'h0; 
  assign _T_1826 = io_in_c_bits_opcode == 3'h5; 
  assign _T_1844 = io_in_c_bits_opcode == 3'h6; 
  assign _T_1859 = io_in_c_bits_size <= 4'h6; 
  assign _T_1867 = _T_1859 & _T_1670; 
  assign _T_1871 = _T_1867 | reset; 
  assign _T_1872 = _T_1871 == 1'h0; 
  assign _T_1941 = _T_1581 ? _T_1859 : 1'h0; 
  assign _T_1958 = _T_1941 | reset; 
  assign _T_1959 = _T_1958 == 1'h0; 
  assign _T_1970 = io_in_c_bits_param <= 3'h2; 
  assign _T_1972 = _T_1970 | reset; 
  assign _T_1973 = _T_1972 == 1'h0; 
  assign _T_1978 = io_in_c_bits_opcode == 3'h7; 
  assign _T_2108 = io_in_c_bits_opcode == 3'h0; 
  assign _T_2118 = io_in_c_bits_param == 3'h0; 
  assign _T_2120 = _T_2118 | reset; 
  assign _T_2121 = _T_2120 == 1'h0; 
  assign _T_2126 = io_in_c_bits_opcode == 3'h1; 
  assign _T_2140 = io_in_c_bits_opcode == 3'h2; 
  assign _T_2158 = io_in_e_bits_sink < 1'h1; 
  assign _T_2160 = _T_2158 | reset; 
  assign _T_2161 = _T_2160 == 1'h0; 
  assign _T_2162 = io_in_a_ready & io_in_a_valid; 
  assign _T_2167 = _T_80[7:3]; 
  assign _T_2168 = io_in_a_bits_opcode[2]; 
  assign _T_2169 = _T_2168 == 1'h0; 
  assign _T_2173 = _T_2171 - 5'h1; 
  assign _T_2174 = _T_2171 == 5'h0; 
  assign _T_2187 = _T_2174 == 1'h0; 
  assign _T_2188 = io_in_a_valid & _T_2187; 
  assign _T_2189 = io_in_a_bits_opcode == _T_2182; 
  assign _T_2191 = _T_2189 | reset; 
  assign _T_2192 = _T_2191 == 1'h0; 
  assign _T_2193 = io_in_a_bits_param == _T_2183; 
  assign _T_2195 = _T_2193 | reset; 
  assign _T_2196 = _T_2195 == 1'h0; 
  assign _T_2197 = io_in_a_bits_size == _T_2184; 
  assign _T_2199 = _T_2197 | reset; 
  assign _T_2200 = _T_2199 == 1'h0; 
  assign _T_2201 = io_in_a_bits_source == _T_2185; 
  assign _T_2203 = _T_2201 | reset; 
  assign _T_2204 = _T_2203 == 1'h0; 
  assign _T_2205 = io_in_a_bits_address == _T_2186; 
  assign _T_2207 = _T_2205 | reset; 
  assign _T_2208 = _T_2207 == 1'h0; 
  assign _T_2210 = _T_2162 & _T_2174; 
  assign _T_2211 = io_in_d_ready & io_in_d_valid; 
  assign _T_2213 = 23'hff << io_in_d_bits_size; 
  assign _T_2214 = _T_2213[7:0]; 
  assign _T_2215 = ~ _T_2214; 
  assign _T_2216 = _T_2215[7:3]; 
  assign _T_2217 = io_in_d_bits_opcode[0]; 
  assign _T_2221 = _T_2219 - 5'h1; 
  assign _T_2222 = _T_2219 == 5'h0; 
  assign _T_2236 = _T_2222 == 1'h0; 
  assign _T_2237 = io_in_d_valid & _T_2236; 
  assign _T_2238 = io_in_d_bits_opcode == _T_2230; 
  assign _T_2240 = _T_2238 | reset; 
  assign _T_2241 = _T_2240 == 1'h0; 
  assign _T_2242 = io_in_d_bits_param == _T_2231; 
  assign _T_2244 = _T_2242 | reset; 
  assign _T_2245 = _T_2244 == 1'h0; 
  assign _T_2246 = io_in_d_bits_size == _T_2232; 
  assign _T_2248 = _T_2246 | reset; 
  assign _T_2249 = _T_2248 == 1'h0; 
  assign _T_2250 = io_in_d_bits_source == _T_2233; 
  assign _T_2252 = _T_2250 | reset; 
  assign _T_2253 = _T_2252 == 1'h0; 
  assign _T_2254 = io_in_d_bits_sink == _T_2234; 
  assign _T_2256 = _T_2254 | reset; 
  assign _T_2257 = _T_2256 == 1'h0; 
  assign _T_2258 = io_in_d_bits_denied == _T_2235; 
  assign _T_2260 = _T_2258 | reset; 
  assign _T_2261 = _T_2260 == 1'h0; 
  assign _T_2263 = _T_2211 & _T_2222; 
  assign _T_2313 = io_in_c_ready & io_in_c_valid; 
  assign _T_2318 = _T_1653[7:3]; 
  assign _T_2319 = io_in_c_bits_opcode[0]; 
  assign _T_2323 = _T_2321 - 5'h1; 
  assign _T_2324 = _T_2321 == 5'h0; 
  assign _T_2337 = _T_2324 == 1'h0; 
  assign _T_2338 = io_in_c_valid & _T_2337; 
  assign _T_2339 = io_in_c_bits_opcode == _T_2332; 
  assign _T_2341 = _T_2339 | reset; 
  assign _T_2342 = _T_2341 == 1'h0; 
  assign _T_2343 = io_in_c_bits_param == _T_2333; 
  assign _T_2345 = _T_2343 | reset; 
  assign _T_2346 = _T_2345 == 1'h0; 
  assign _T_2347 = io_in_c_bits_size == _T_2334; 
  assign _T_2349 = _T_2347 | reset; 
  assign _T_2350 = _T_2349 == 1'h0; 
  assign _T_2351 = io_in_c_bits_source == _T_2335; 
  assign _T_2353 = _T_2351 | reset; 
  assign _T_2354 = _T_2353 == 1'h0; 
  assign _T_2355 = io_in_c_bits_address == _T_2336; 
  assign _T_2357 = _T_2355 | reset; 
  assign _T_2358 = _T_2357 == 1'h0; 
  assign _T_2360 = _T_2313 & _T_2324; 
  assign _T_2373 = _T_2371 - 5'h1; 
  assign _T_2374 = _T_2371 == 5'h0; 
  assign _T_2392 = _T_2390 - 5'h1; 
  assign _T_2393 = _T_2390 == 5'h0; 
  assign _T_2403 = _T_2162 & _T_2374; 
  assign _T_2405 = 128'h1 << io_in_a_bits_source; 
  assign _T_2406 = _T_2361 >> io_in_a_bits_source; 
  assign _T_2407 = _T_2406[0]; 
  assign _T_2408 = _T_2407 == 1'h0; 
  assign _T_2410 = _T_2408 | reset; 
  assign _T_2411 = _T_2410 == 1'h0; 
  assign _GEN_27 = _T_2403 ? _T_2405 : 128'h0; 
  assign _T_2415 = _T_2211 & _T_2393; 
  assign _T_2417 = _T_900 == 1'h0; 
  assign _T_2418 = _T_2415 & _T_2417; 
  assign _T_2419 = 128'h1 << io_in_d_bits_source; 
  assign _T_2420 = _GEN_27 | _T_2361; 
  assign _T_2421 = _T_2420 >> io_in_d_bits_source; 
  assign _T_2422 = _T_2421[0]; 
  assign _T_2424 = _T_2422 | reset; 
  assign _T_2425 = _T_2424 == 1'h0; 
  assign _GEN_28 = _T_2418 ? _T_2419 : 128'h0; 
  assign _T_2426 = _GEN_27 != _GEN_28; 
  assign _T_2427 = _GEN_27 != 128'h0; 
  assign _T_2428 = _T_2427 == 1'h0; 
  assign _T_2429 = _T_2426 | _T_2428; 
  assign _T_2431 = _T_2429 | reset; 
  assign _T_2432 = _T_2431 == 1'h0; 
  assign _T_2433 = _T_2361 | _GEN_27; 
  assign _T_2434 = ~ _GEN_28; 
  assign _T_2435 = _T_2433 & _T_2434; 
  assign _T_2437 = _T_2361 != 128'h0; 
  assign _T_2438 = _T_2437 == 1'h0; 
  assign _T_2439 = plusarg_reader_out == 32'h0; 
  assign _T_2440 = _T_2438 | _T_2439; 
  assign _T_2441 = _T_2436 < plusarg_reader_out; 
  assign _T_2442 = _T_2440 | _T_2441; 
  assign _T_2444 = _T_2442 | reset; 
  assign _T_2445 = _T_2444 == 1'h0; 
  assign _T_2447 = _T_2436 + 32'h1; 
  assign _T_2450 = _T_2162 | _T_2211; 
  assign _T_2462 = _T_2460 - 5'h1; 
  assign _T_2463 = _T_2460 == 5'h0; 
  assign _T_2473 = _T_2211 & _T_2463; 
  assign _T_2474 = io_in_d_bits_opcode[2]; 
  assign _T_2475 = io_in_d_bits_opcode[1]; 
  assign _T_2476 = _T_2475 == 1'h0; 
  assign _T_2477 = _T_2474 & _T_2476; 
  assign _T_2478 = _T_2473 & _T_2477; 
  assign _T_2479 = 2'h1 << io_in_d_bits_sink; 
  assign _T_2480 = _T_2451 >> io_in_d_bits_sink; 
  assign _T_2482 = _T_2480 == 1'h0; 
  assign _T_2484 = _T_2482 | reset; 
  assign _T_2485 = _T_2484 == 1'h0; 
  assign _GEN_31 = _T_2478 ? _T_2479 : 2'h0; 
  assign _T_2487 = io_in_e_ready & io_in_e_valid; 
  assign _T_2490 = 2'h1 << io_in_e_bits_sink; 
  assign _T_2471 = _GEN_31[0]; 
  assign _T_2491 = _T_2471 | _T_2451; 
  assign _T_2492 = _T_2491 >> io_in_e_bits_sink; 
  assign _T_2495 = _T_2492 | reset; 
  assign _T_2496 = _T_2495 == 1'h0; 
  assign _GEN_32 = _T_2487 ? _T_2490 : 2'h0; 
  assign _T_2497 = _T_2451 | _T_2471; 
  assign _T_2486 = _GEN_32[0]; 
  assign _T_2498 = ~ _T_2486; 
  assign _T_2499 = _T_2497 & _T_2498; 
  assign _GEN_35 = io_in_a_valid & _T_277; 
  assign _GEN_49 = io_in_a_valid & _T_416; 
  assign _GEN_65 = io_in_a_valid & _T_559; 
  assign _GEN_75 = io_in_a_valid & _T_604; 
  assign _GEN_85 = io_in_a_valid & _T_650; 
  assign _GEN_95 = io_in_a_valid & _T_698; 
  assign _GEN_105 = io_in_a_valid & _T_739; 
  assign _GEN_115 = io_in_a_valid & _T_780; 
  assign _GEN_123 = io_in_d_valid & _T_900; 
  assign _GEN_133 = io_in_d_valid & _T_920; 
  assign _GEN_145 = io_in_d_valid & _T_948; 
  assign _GEN_157 = io_in_d_valid & _T_977; 
  assign _GEN_163 = io_in_d_valid & _T_994; 
  assign _GEN_169 = io_in_d_valid & _T_1012; 
  assign _GEN_175 = io_in_c_valid & _T_1804; 
  assign _GEN_187 = io_in_c_valid & _T_1826; 
  assign _GEN_197 = io_in_c_valid & _T_1844; 
  assign _GEN_211 = io_in_c_valid & _T_1978; 
  assign _GEN_223 = io_in_c_valid & _T_2108; 
  assign _GEN_233 = io_in_c_valid & _T_2126; 
  assign _GEN_241 = io_in_c_valid & _T_2140; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2171 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_2182 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2183 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_2184 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_2185 = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_2186 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_2219 = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_2230 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_2231 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_2232 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_2233 = _RAND_10[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_2234 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_2235 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_2321 = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_2332 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_2333 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_2334 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_2335 = _RAND_17[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_2336 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {4{`RANDOM}};
  _T_2361 = _RAND_19[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_2371 = _RAND_20[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_2390 = _RAND_21[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_2436 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_2451 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_2460 = _RAND_24[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_2171 <= 5'h0;
    end else begin
      if (_T_2162) begin
        if (_T_2174) begin
          if (_T_2169) begin
            _T_2171 <= _T_2167;
          end else begin
            _T_2171 <= 5'h0;
          end
        end else begin
          _T_2171 <= _T_2173;
        end
      end
    end
    if (_T_2210) begin
      _T_2182 <= io_in_a_bits_opcode;
    end
    if (_T_2210) begin
      _T_2183 <= io_in_a_bits_param;
    end
    if (_T_2210) begin
      _T_2184 <= io_in_a_bits_size;
    end
    if (_T_2210) begin
      _T_2185 <= io_in_a_bits_source;
    end
    if (_T_2210) begin
      _T_2186 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_2219 <= 5'h0;
    end else begin
      if (_T_2211) begin
        if (_T_2222) begin
          if (_T_2217) begin
            _T_2219 <= _T_2216;
          end else begin
            _T_2219 <= 5'h0;
          end
        end else begin
          _T_2219 <= _T_2221;
        end
      end
    end
    if (_T_2263) begin
      _T_2230 <= io_in_d_bits_opcode;
    end
    if (_T_2263) begin
      _T_2231 <= io_in_d_bits_param;
    end
    if (_T_2263) begin
      _T_2232 <= io_in_d_bits_size;
    end
    if (_T_2263) begin
      _T_2233 <= io_in_d_bits_source;
    end
    if (_T_2263) begin
      _T_2234 <= io_in_d_bits_sink;
    end
    if (_T_2263) begin
      _T_2235 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_2321 <= 5'h0;
    end else begin
      if (_T_2313) begin
        if (_T_2324) begin
          if (_T_2319) begin
            _T_2321 <= _T_2318;
          end else begin
            _T_2321 <= 5'h0;
          end
        end else begin
          _T_2321 <= _T_2323;
        end
      end
    end
    if (_T_2360) begin
      _T_2332 <= io_in_c_bits_opcode;
    end
    if (_T_2360) begin
      _T_2333 <= io_in_c_bits_param;
    end
    if (_T_2360) begin
      _T_2334 <= io_in_c_bits_size;
    end
    if (_T_2360) begin
      _T_2335 <= io_in_c_bits_source;
    end
    if (_T_2360) begin
      _T_2336 <= io_in_c_bits_address;
    end
    if (reset) begin
      _T_2361 <= 128'h0;
    end else begin
      _T_2361 <= _T_2435;
    end
    if (reset) begin
      _T_2371 <= 5'h0;
    end else begin
      if (_T_2162) begin
        if (_T_2374) begin
          if (_T_2169) begin
            _T_2371 <= _T_2167;
          end else begin
            _T_2371 <= 5'h0;
          end
        end else begin
          _T_2371 <= _T_2373;
        end
      end
    end
    if (reset) begin
      _T_2390 <= 5'h0;
    end else begin
      if (_T_2211) begin
        if (_T_2393) begin
          if (_T_2217) begin
            _T_2390 <= _T_2216;
          end else begin
            _T_2390 <= 5'h0;
          end
        end else begin
          _T_2390 <= _T_2392;
        end
      end
    end
    if (reset) begin
      _T_2436 <= 32'h0;
    end else begin
      if (_T_2450) begin
        _T_2436 <= 32'h0;
      end else begin
        _T_2436 <= _T_2447;
      end
    end
    if (reset) begin
      _T_2451 <= 1'h0;
    end else begin
      _T_2451 <= _T_2499;
    end
    if (reset) begin
      _T_2460 <= 5'h0;
    end else begin
      if (_T_2211) begin
        if (_T_2463) begin
          if (_T_2217) begin
            _T_2460 <= _T_2216;
          end else begin
            _T_2460 <= 5'h0;
          end
        end else begin
          _T_2460 <= _T_2462;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel has invalid opcode (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:39 assert (TLMessages.isA(bundle.opcode), \"'A' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:46 assert (visible(edge.address(bundle), bundle.source, edge), \"'A' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_305) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_305) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_392) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_392) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_399) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_399) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_406) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_406) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_411) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_411) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:56 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_305) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_305) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_392) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_392) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_399) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_399) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_406) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_406) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_549) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_549) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_411) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_411) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:68 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_585) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_585) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_595) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_595) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_599) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:77 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_635) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_635) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_595) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_595) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_599) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_635) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_635) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_595) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_595) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_697) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_697) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_724) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_724) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_734) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_734) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_599) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_724) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_724) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_775) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_775) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_599) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_305) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_305) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_599) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:117 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_826) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_826) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_903) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_903) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_907) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_907) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_911) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_911) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_915) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_915) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_919) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_919) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_903) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_903) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_926) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:285 assert (sink_ok, \"'D' channel Grant carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_926) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_907) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_907) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_934) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_934) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_938) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_938) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_915) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_915) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is denied (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:290 assert (deny_put_ok || !bundle.denied, \"'D' channel Grant is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_903) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_903) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_926) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:295 assert (sink_ok, \"'D' channel GrantData carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_926) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_907) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_907) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_934) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_934) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_938) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_938) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_971) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_971) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:300 assert (deny_get_ok || !bundle.denied, \"'D' channel GrantData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_157 & _T_903) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_157 & _T_903) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_157 & _T_911) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_157 & _T_911) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_157 & _T_915) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_157 & _T_915) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is denied (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:308 assert (deny_put_ok || !bundle.denied, \"'D' channel AccessAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_903) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_903) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_911) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_911) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_971) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_971) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:316 assert (deny_get_ok || !bundle.denied, \"'D' channel AccessAckData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_169 & _T_903) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_169 & _T_903) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_169 & _T_911) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_169 & _T_911) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_169 & _T_915) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_169 & _T_915) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is denied (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:324 assert (deny_put_ok || !bundle.denied, \"'D' channel HintAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel has invalid opcode (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:122 assert (TLMessages.isB(bundle.opcode), \"'B' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:124 assert (visible(edge.address(bundle), bundle.source, edge), \"'B' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Probe type unsupported by client (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:133 assert (edge.client.supportsProbe(bundle.source, bundle.size), \"'B' channel carries Probe type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:134 assert (address_ok, \"'B' channel Probe carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries source that is not first source (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:135 assert (legal_source, \"'B' channel Probe carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:136 assert (is_aligned, \"'B' channel Probe address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:137 assert (TLPermissions.isCap(bundle.param), \"'B' channel Probe carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe contains invalid mask (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:138 assert (bundle.mask === mask, \"'B' channel Probe contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe is corrupt (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:139 assert (!bundle.corrupt, \"'B' channel Probe is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Get type unsupported by client (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:143 assert (edge.client.supportsGet(bundle.source, bundle.size), \"'B' channel carries Get type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries unmanaged address (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:144 assert (address_ok, \"'B' channel Get carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries source that is not first source (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:145 assert (legal_source, \"'B' channel Get carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:146 assert (is_aligned, \"'B' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries invalid param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:147 assert (bundle.param === UInt(0), \"'B' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get contains invalid mask (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:148 assert (bundle.mask === mask, \"'B' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get is corrupt (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:149 assert (!bundle.corrupt, \"'B' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutFull type unsupported by client (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:153 assert (edge.client.supportsPutFull(bundle.source, bundle.size), \"'B' channel carries PutFull type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries unmanaged address (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:154 assert (address_ok, \"'B' channel PutFull carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries source that is not first source (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:155 assert (legal_source, \"'B' channel PutFull carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:156 assert (is_aligned, \"'B' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries invalid param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:157 assert (bundle.param === UInt(0), \"'B' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull contains invalid mask (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:158 assert (bundle.mask === mask, \"'B' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutPartial type unsupported by client (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:162 assert (edge.client.supportsPutPartial(bundle.source, bundle.size), \"'B' channel carries PutPartial type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:163 assert (address_ok, \"'B' channel PutPartial carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:164 assert (legal_source, \"'B' channel PutPartial carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:165 assert (is_aligned, \"'B' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries invalid param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:166 assert (bundle.param === UInt(0), \"'B' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial contains invalid mask (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:167 assert ((bundle.mask & ~mask) === UInt(0), \"'B' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Arithmetic type unsupported by client (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:171 assert (edge.client.supportsArithmetic(bundle.source, bundle.size), \"'B' channel carries Arithmetic type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:172 assert (address_ok, \"'B' channel Arithmetic carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:173 assert (legal_source, \"'B' channel Arithmetic carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:174 assert (is_aligned, \"'B' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries invalid opcode param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:175 assert (TLAtomics.isArithmetic(bundle.param), \"'B' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:176 assert (bundle.mask === mask, \"'B' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Logical type unsupported by client (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:180 assert (edge.client.supportsLogical(bundle.source, bundle.size), \"'B' channel carries Logical type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries unmanaged address (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:181 assert (address_ok, \"'B' channel Logical carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries source that is not first source (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:182 assert (legal_source, \"'B' channel Logical carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:183 assert (is_aligned, \"'B' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries invalid opcode param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:184 assert (TLAtomics.isLogical(bundle.param), \"'B' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical contains invalid mask (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:185 assert (bundle.mask === mask, \"'B' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Hint type unsupported by client (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:189 assert (edge.client.supportsHint(bundle.source, bundle.size), \"'B' channel carries Hint type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries unmanaged address (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:190 assert (address_ok, \"'B' channel Hint carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries source that is not first source (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:191 assert (legal_source, \"'B' channel Hint carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:192 assert (is_aligned, \"'B' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint contains invalid mask (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:193 assert (bundle.mask === mask, \"'B' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint is corrupt (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:194 assert (!bundle.corrupt, \"'B' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel has invalid opcode (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:199 assert (TLMessages.isC(bundle.opcode), \"'C' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:205 assert (visible(edge.address(bundle), bundle.source, edge), \"'C' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1807) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:208 assert (address_ok, \"'C' channel ProbeAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1807) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1810) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:209 assert (source_ok, \"'C' channel ProbeAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1810) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1814) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:210 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1814) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1817) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:211 assert (is_aligned, \"'C' channel ProbeAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1817) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1821) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:212 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAck carries invalid report param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1821) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1825) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck is corrupt (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:213 assert (!bundle.corrupt, \"'C' channel ProbeAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1825) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_187 & _T_1807) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:217 assert (address_ok, \"'C' channel ProbeAckData carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_187 & _T_1807) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_187 & _T_1810) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:218 assert (source_ok, \"'C' channel ProbeAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_187 & _T_1810) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_187 & _T_1814) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:219 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAckData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_187 & _T_1814) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_187 & _T_1817) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:220 assert (is_aligned, \"'C' channel ProbeAckData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_187 & _T_1817) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_187 & _T_1821) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:221 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAckData carries invalid report param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_187 & _T_1821) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1872) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:225 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries Release type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1872) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1959) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:226 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1959) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1810) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:227 assert (source_ok, \"'C' channel Release carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1810) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1814) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:228 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel Release smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1814) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1817) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:229 assert (is_aligned, \"'C' channel Release address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1817) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1973) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid shrink param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:230 assert (TLPermissions.isShrink(bundle.param), \"'C' channel Release carries invalid shrink param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1973) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1825) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release is corrupt (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:231 assert (!bundle.corrupt, \"'C' channel Release is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1825) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1872) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:235 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries ReleaseData type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1872) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1959) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:236 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1959) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1810) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:237 assert (source_ok, \"'C' channel ReleaseData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1810) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1814) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:238 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ReleaseData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1814) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1817) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:239 assert (is_aligned, \"'C' channel ReleaseData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1817) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1973) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid shrink param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:240 assert (TLPermissions.isShrink(bundle.param), \"'C' channel ReleaseData carries invalid shrink param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1973) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_1807) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:244 assert (address_ok, \"'C' channel AccessAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_1807) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_1810) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:245 assert (source_ok, \"'C' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_1810) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_1817) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:246 assert (is_aligned, \"'C' channel AccessAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_1817) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_2121) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:247 assert (bundle.param === UInt(0), \"'C' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_2121) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_1825) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck is corrupt (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:248 assert (!bundle.corrupt, \"'C' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_1825) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_1807) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:252 assert (address_ok, \"'C' channel AccessAckData carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_1807) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_1810) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:253 assert (source_ok, \"'C' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_1810) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_1817) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:254 assert (is_aligned, \"'C' channel AccessAckData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_1817) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_2121) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:255 assert (bundle.param === UInt(0), \"'C' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_2121) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1807) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:259 assert (address_ok, \"'C' channel HintAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1807) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1810) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:260 assert (source_ok, \"'C' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1810) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1817) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:261 assert (is_aligned, \"'C' channel HintAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1817) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_2121) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:262 assert (bundle.param === UInt(0), \"'C' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_2121) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1825) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck is corrupt (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:263 assert (!bundle.corrupt, \"'C' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1825) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_e_valid & _T_2161) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channels carries invalid sink ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:330 assert (sink_ok, \"'E' channels carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_e_valid & _T_2161) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2188 & _T_2192) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2188 & _T_2192) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2188 & _T_2196) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2188 & _T_2196) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2188 & _T_2200) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2188 & _T_2200) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2188 & _T_2204) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2188 & _T_2204) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2188 & _T_2208) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2188 & _T_2208) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2237 & _T_2241) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2237 & _T_2241) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2237 & _T_2245) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2237 & _T_2245) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2237 & _T_2249) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2237 & _T_2249) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2237 & _T_2253) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2237 & _T_2253) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2237 & _T_2257) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2237 & _T_2257) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2237 & _T_2261) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2237 & _T_2261) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:378 assert (b.bits.opcode === opcode, \"'B' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:379 assert (b.bits.param  === param,  \"'B' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel size changed within multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:380 assert (b.bits.size   === size,   \"'B' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel source changed within multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:381 assert (b.bits.source === source, \"'B' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:382 assert (b.bits.address=== address,\"'B' channel addresss changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2338 & _T_2342) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:401 assert (c.bits.opcode === opcode, \"'C' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2338 & _T_2342) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2338 & _T_2346) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:402 assert (c.bits.param  === param,  \"'C' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2338 & _T_2346) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2338 & _T_2350) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:403 assert (c.bits.size   === size,   \"'C' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2338 & _T_2350) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2338 & _T_2354) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:404 assert (c.bits.source === source, \"'C' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2338 & _T_2354) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2338 & _T_2358) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:405 assert (c.bits.address=== address,\"'C' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2338 & _T_2358) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2403 & _T_2411) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2403 & _T_2411) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2418 & _T_2425) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2418 & _T_2425) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2432) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2432) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2445) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:479 assert (!inflight.orR || limit === UInt(0) || watchdog < limit, \"TileLink timeout expired\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2445) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2478 & _T_2485) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:494 assert(!inflight(bundle.d.bits.sink), \"'D' channel re-used a sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2478 & _T_2485) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2487 & _T_2496) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at ChiplinkTest.scala:362:79)\n    at Monitor.scala:500 assert((d_set | inflight)(bundle.e.bits.sink), \"'E' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2487 & _T_2496) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLMonitor_16( 
  input         clock, 
  input         reset, 
  input         io_in_a_ready, 
  input         io_in_a_valid, 
  input  [2:0]  io_in_a_bits_opcode, 
  input  [2:0]  io_in_a_bits_param, 
  input  [3:0]  io_in_a_bits_size, 
  input  [5:0]  io_in_a_bits_source, 
  input  [31:0] io_in_a_bits_address, 
  input  [7:0]  io_in_a_bits_mask, 
  input         io_in_c_ready, 
  input         io_in_c_valid, 
  input  [2:0]  io_in_c_bits_opcode, 
  input  [2:0]  io_in_c_bits_param, 
  input  [3:0]  io_in_c_bits_size, 
  input  [5:0]  io_in_c_bits_source, 
  input  [31:0] io_in_c_bits_address, 
  input         io_in_c_bits_corrupt, 
  input         io_in_d_ready, 
  input         io_in_d_valid, 
  input  [2:0]  io_in_d_bits_opcode, 
  input  [1:0]  io_in_d_bits_param, 
  input  [3:0]  io_in_d_bits_size, 
  input  [5:0]  io_in_d_bits_source, 
  input         io_in_d_bits_sink, 
  input         io_in_d_bits_denied, 
  input         io_in_d_bits_corrupt, 
  input         io_in_e_ready, 
  input         io_in_e_valid, 
  input         io_in_e_bits_sink 
);
  wire [31:0] plusarg_reader_out; 
  wire [2:0] _T_7; 
  wire  _T_8; 
  wire  _T_16; 
  wire  _T_24; 
  wire  _T_32; 
  wire  _T_40; 
  wire  _T_48; 
  wire  _T_56; 
  wire  _T_64; 
  wire  _T_70; 
  wire  _T_71; 
  wire  _T_72; 
  wire  _T_73; 
  wire  _T_74; 
  wire  _T_75; 
  wire  _T_76; 
  wire [22:0] _T_78; 
  wire [7:0] _T_79; 
  wire [7:0] _T_80; 
  wire [31:0] _GEN_33; 
  wire [31:0] _T_81; 
  wire  _T_82; 
  wire [1:0] _T_84; 
  wire [3:0] _T_85; 
  wire [2:0] _T_86; 
  wire [2:0] _T_87; 
  wire  _T_88; 
  wire  _T_89; 
  wire  _T_90; 
  wire  _T_91; 
  wire  _T_93; 
  wire  _T_94; 
  wire  _T_96; 
  wire  _T_97; 
  wire  _T_98; 
  wire  _T_99; 
  wire  _T_100; 
  wire  _T_101; 
  wire  _T_102; 
  wire  _T_103; 
  wire  _T_104; 
  wire  _T_105; 
  wire  _T_106; 
  wire  _T_107; 
  wire  _T_108; 
  wire  _T_109; 
  wire  _T_110; 
  wire  _T_111; 
  wire  _T_112; 
  wire  _T_113; 
  wire  _T_114; 
  wire  _T_115; 
  wire  _T_116; 
  wire  _T_117; 
  wire  _T_118; 
  wire  _T_119; 
  wire  _T_120; 
  wire  _T_121; 
  wire  _T_122; 
  wire  _T_123; 
  wire  _T_124; 
  wire  _T_125; 
  wire  _T_126; 
  wire  _T_127; 
  wire  _T_128; 
  wire  _T_129; 
  wire  _T_130; 
  wire  _T_131; 
  wire  _T_132; 
  wire  _T_133; 
  wire  _T_134; 
  wire  _T_135; 
  wire  _T_136; 
  wire  _T_137; 
  wire  _T_138; 
  wire  _T_139; 
  wire [7:0] _T_146; 
  wire  _T_277; 
  wire [31:0] _T_279; 
  wire [32:0] _T_280; 
  wire [32:0] _T_281; 
  wire [32:0] _T_282; 
  wire  _T_283; 
  wire [31:0] _T_284; 
  wire [32:0] _T_285; 
  wire [32:0] _T_286; 
  wire [32:0] _T_287; 
  wire  _T_288; 
  wire  _T_289; 
  wire  _T_292; 
  wire [31:0] _T_295; 
  wire [32:0] _T_296; 
  wire [32:0] _T_297; 
  wire [32:0] _T_298; 
  wire  _T_299; 
  wire  _T_300; 
  wire  _T_304; 
  wire  _T_305; 
  wire  _T_374; 
  wire  _T_391; 
  wire  _T_392; 
  wire  _T_394; 
  wire  _T_395; 
  wire  _T_398; 
  wire  _T_399; 
  wire  _T_401; 
  wire  _T_402; 
  wire  _T_403; 
  wire  _T_405; 
  wire  _T_406; 
  wire [7:0] _T_407; 
  wire  _T_408; 
  wire  _T_410; 
  wire  _T_411; 
  wire  _T_416; 
  wire  _T_546; 
  wire  _T_548; 
  wire  _T_549; 
  wire  _T_559; 
  wire  _T_580; 
  wire  _T_581; 
  wire  _T_584; 
  wire  _T_585; 
  wire  _T_592; 
  wire  _T_594; 
  wire  _T_595; 
  wire  _T_596; 
  wire  _T_598; 
  wire  _T_599; 
  wire  _T_604; 
  wire  _T_619; 
  wire  _T_620; 
  wire  _T_622; 
  wire  _T_630; 
  wire  _T_632; 
  wire  _T_634; 
  wire  _T_635; 
  wire  _T_650; 
  wire [7:0] _T_692; 
  wire [7:0] _T_693; 
  wire  _T_694; 
  wire  _T_696; 
  wire  _T_697; 
  wire  _T_698; 
  wire  _T_700; 
  wire  _T_720; 
  wire  _T_723; 
  wire  _T_724; 
  wire  _T_731; 
  wire  _T_733; 
  wire  _T_734; 
  wire  _T_739; 
  wire  _T_772; 
  wire  _T_774; 
  wire  _T_775; 
  wire  _T_780; 
  wire  _T_826; 
  wire  _T_828; 
  wire  _T_829; 
  wire [2:0] _T_832; 
  wire  _T_833; 
  wire  _T_841; 
  wire  _T_849; 
  wire  _T_857; 
  wire  _T_865; 
  wire  _T_873; 
  wire  _T_881; 
  wire  _T_889; 
  wire  _T_895; 
  wire  _T_896; 
  wire  _T_897; 
  wire  _T_898; 
  wire  _T_899; 
  wire  _T_900; 
  wire  _T_901; 
  wire  _T_902; 
  wire  _T_903; 
  wire  _T_905; 
  wire  _T_906; 
  wire  _T_907; 
  wire  _T_909; 
  wire  _T_910; 
  wire  _T_911; 
  wire  _T_913; 
  wire  _T_914; 
  wire  _T_915; 
  wire  _T_917; 
  wire  _T_918; 
  wire  _T_919; 
  wire  _T_921; 
  wire  _T_922; 
  wire  _T_923; 
  wire  _T_928; 
  wire  _T_929; 
  wire  _T_934; 
  wire  _T_936; 
  wire  _T_937; 
  wire  _T_938; 
  wire  _T_940; 
  wire  _T_941; 
  wire  _T_951; 
  wire  _T_971; 
  wire  _T_973; 
  wire  _T_974; 
  wire  _T_980; 
  wire  _T_997; 
  wire  _T_1015; 
  wire [2:0] _T_1583; 
  wire  _T_1584; 
  wire  _T_1592; 
  wire  _T_1600; 
  wire  _T_1608; 
  wire  _T_1616; 
  wire  _T_1624; 
  wire  _T_1632; 
  wire  _T_1640; 
  wire  _T_1646; 
  wire  _T_1647; 
  wire  _T_1648; 
  wire  _T_1649; 
  wire  _T_1650; 
  wire  _T_1651; 
  wire  _T_1652; 
  wire [22:0] _T_1654; 
  wire [7:0] _T_1655; 
  wire [7:0] _T_1656; 
  wire [31:0] _GEN_34; 
  wire [31:0] _T_1657; 
  wire  _T_1658; 
  wire [31:0] _T_1659; 
  wire [32:0] _T_1660; 
  wire [32:0] _T_1661; 
  wire [32:0] _T_1662; 
  wire  _T_1663; 
  wire [31:0] _T_1664; 
  wire [32:0] _T_1665; 
  wire [32:0] _T_1666; 
  wire [32:0] _T_1667; 
  wire  _T_1668; 
  wire [31:0] _T_1669; 
  wire [32:0] _T_1670; 
  wire [32:0] _T_1671; 
  wire [32:0] _T_1672; 
  wire  _T_1673; 
  wire  _T_1675; 
  wire  _T_1676; 
  wire  _T_1807; 
  wire  _T_1809; 
  wire  _T_1810; 
  wire  _T_1812; 
  wire  _T_1813; 
  wire  _T_1814; 
  wire  _T_1816; 
  wire  _T_1817; 
  wire  _T_1819; 
  wire  _T_1820; 
  wire  _T_1821; 
  wire  _T_1823; 
  wire  _T_1824; 
  wire  _T_1825; 
  wire  _T_1827; 
  wire  _T_1828; 
  wire  _T_1829; 
  wire  _T_1847; 
  wire  _T_1862; 
  wire  _T_1870; 
  wire  _T_1874; 
  wire  _T_1875; 
  wire  _T_1944; 
  wire  _T_1961; 
  wire  _T_1962; 
  wire  _T_1973; 
  wire  _T_1975; 
  wire  _T_1976; 
  wire  _T_1981; 
  wire  _T_2111; 
  wire  _T_2121; 
  wire  _T_2123; 
  wire  _T_2124; 
  wire  _T_2129; 
  wire  _T_2143; 
  wire  _T_2161; 
  wire  _T_2163; 
  wire  _T_2164; 
  wire  _T_2165; 
  wire [4:0] _T_2170; 
  wire  _T_2171; 
  wire  _T_2172; 
  reg [4:0] _T_2174; 
  reg [31:0] _RAND_0;
  wire [4:0] _T_2176; 
  wire  _T_2177; 
  reg [2:0] _T_2185; 
  reg [31:0] _RAND_1;
  reg [2:0] _T_2186; 
  reg [31:0] _RAND_2;
  reg [3:0] _T_2187; 
  reg [31:0] _RAND_3;
  reg [5:0] _T_2188; 
  reg [31:0] _RAND_4;
  reg [31:0] _T_2189; 
  reg [31:0] _RAND_5;
  wire  _T_2190; 
  wire  _T_2191; 
  wire  _T_2192; 
  wire  _T_2194; 
  wire  _T_2195; 
  wire  _T_2196; 
  wire  _T_2198; 
  wire  _T_2199; 
  wire  _T_2200; 
  wire  _T_2202; 
  wire  _T_2203; 
  wire  _T_2204; 
  wire  _T_2206; 
  wire  _T_2207; 
  wire  _T_2208; 
  wire  _T_2210; 
  wire  _T_2211; 
  wire  _T_2213; 
  wire  _T_2214; 
  wire [22:0] _T_2216; 
  wire [7:0] _T_2217; 
  wire [7:0] _T_2218; 
  wire [4:0] _T_2219; 
  wire  _T_2220; 
  reg [4:0] _T_2222; 
  reg [31:0] _RAND_6;
  wire [4:0] _T_2224; 
  wire  _T_2225; 
  reg [2:0] _T_2233; 
  reg [31:0] _RAND_7;
  reg [1:0] _T_2234; 
  reg [31:0] _RAND_8;
  reg [3:0] _T_2235; 
  reg [31:0] _RAND_9;
  reg [5:0] _T_2236; 
  reg [31:0] _RAND_10;
  reg  _T_2237; 
  reg [31:0] _RAND_11;
  reg  _T_2238; 
  reg [31:0] _RAND_12;
  wire  _T_2239; 
  wire  _T_2240; 
  wire  _T_2241; 
  wire  _T_2243; 
  wire  _T_2244; 
  wire  _T_2245; 
  wire  _T_2247; 
  wire  _T_2248; 
  wire  _T_2249; 
  wire  _T_2251; 
  wire  _T_2252; 
  wire  _T_2253; 
  wire  _T_2255; 
  wire  _T_2256; 
  wire  _T_2257; 
  wire  _T_2259; 
  wire  _T_2260; 
  wire  _T_2261; 
  wire  _T_2263; 
  wire  _T_2264; 
  wire  _T_2266; 
  wire  _T_2316; 
  wire [4:0] _T_2321; 
  wire  _T_2322; 
  reg [4:0] _T_2324; 
  reg [31:0] _RAND_13;
  wire [4:0] _T_2326; 
  wire  _T_2327; 
  reg [2:0] _T_2335; 
  reg [31:0] _RAND_14;
  reg [2:0] _T_2336; 
  reg [31:0] _RAND_15;
  reg [3:0] _T_2337; 
  reg [31:0] _RAND_16;
  reg [5:0] _T_2338; 
  reg [31:0] _RAND_17;
  reg [31:0] _T_2339; 
  reg [31:0] _RAND_18;
  wire  _T_2340; 
  wire  _T_2341; 
  wire  _T_2342; 
  wire  _T_2344; 
  wire  _T_2345; 
  wire  _T_2346; 
  wire  _T_2348; 
  wire  _T_2349; 
  wire  _T_2350; 
  wire  _T_2352; 
  wire  _T_2353; 
  wire  _T_2354; 
  wire  _T_2356; 
  wire  _T_2357; 
  wire  _T_2358; 
  wire  _T_2360; 
  wire  _T_2361; 
  wire  _T_2363; 
  reg [63:0] _T_2364; 
  reg [63:0] _RAND_19;
  reg [4:0] _T_2374; 
  reg [31:0] _RAND_20;
  wire [4:0] _T_2376; 
  wire  _T_2377; 
  reg [4:0] _T_2393; 
  reg [31:0] _RAND_21;
  wire [4:0] _T_2395; 
  wire  _T_2396; 
  wire  _T_2406; 
  wire [63:0] _T_2408; 
  wire [63:0] _T_2409; 
  wire  _T_2410; 
  wire  _T_2411; 
  wire  _T_2413; 
  wire  _T_2414; 
  wire [63:0] _GEN_27; 
  wire  _T_2418; 
  wire  _T_2420; 
  wire  _T_2421; 
  wire [63:0] _T_2422; 
  wire [63:0] _T_2423; 
  wire [63:0] _T_2424; 
  wire  _T_2425; 
  wire  _T_2427; 
  wire  _T_2428; 
  wire [63:0] _GEN_28; 
  wire  _T_2429; 
  wire  _T_2430; 
  wire  _T_2431; 
  wire  _T_2432; 
  wire  _T_2434; 
  wire  _T_2435; 
  wire [63:0] _T_2436; 
  wire [63:0] _T_2437; 
  wire [63:0] _T_2438; 
  reg [31:0] _T_2439; 
  reg [31:0] _RAND_22;
  wire  _T_2440; 
  wire  _T_2441; 
  wire  _T_2442; 
  wire  _T_2443; 
  wire  _T_2444; 
  wire  _T_2445; 
  wire  _T_2447; 
  wire  _T_2448; 
  wire [31:0] _T_2450; 
  wire  _T_2453; 
  reg  _T_2454; 
  reg [31:0] _RAND_23;
  reg [4:0] _T_2463; 
  reg [31:0] _RAND_24;
  wire [4:0] _T_2465; 
  wire  _T_2466; 
  wire  _T_2476; 
  wire  _T_2477; 
  wire  _T_2478; 
  wire  _T_2479; 
  wire  _T_2480; 
  wire  _T_2481; 
  wire [1:0] _T_2482; 
  wire  _T_2483; 
  wire  _T_2485; 
  wire  _T_2487; 
  wire  _T_2488; 
  wire [1:0] _GEN_31; 
  wire  _T_2490; 
  wire [1:0] _T_2493; 
  wire  _T_2474; 
  wire  _T_2494; 
  wire  _T_2495; 
  wire  _T_2498; 
  wire  _T_2499; 
  wire [1:0] _GEN_32; 
  wire  _T_2500; 
  wire  _T_2489; 
  wire  _T_2501; 
  wire  _T_2502; 
  wire  _GEN_35; 
  wire  _GEN_49; 
  wire  _GEN_65; 
  wire  _GEN_75; 
  wire  _GEN_85; 
  wire  _GEN_95; 
  wire  _GEN_105; 
  wire  _GEN_115; 
  wire  _GEN_123; 
  wire  _GEN_133; 
  wire  _GEN_145; 
  wire  _GEN_157; 
  wire  _GEN_163; 
  wire  _GEN_169; 
  wire  _GEN_175; 
  wire  _GEN_187; 
  wire  _GEN_197; 
  wire  _GEN_211; 
  wire  _GEN_223; 
  wire  _GEN_233; 
  wire  _GEN_241; 
  dual_plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0)) plusarg_reader ( 
    .out(plusarg_reader_out)
  );
  assign _T_7 = io_in_a_bits_source[5:3]; 
  assign _T_8 = _T_7 == 3'h0; 
  assign _T_16 = _T_7 == 3'h1; 
  assign _T_24 = _T_7 == 3'h2; 
  assign _T_32 = _T_7 == 3'h3; 
  assign _T_40 = _T_7 == 3'h4; 
  assign _T_48 = _T_7 == 3'h5; 
  assign _T_56 = _T_7 == 3'h6; 
  assign _T_64 = _T_7 == 3'h7; 
  assign _T_70 = _T_8 | _T_16; 
  assign _T_71 = _T_70 | _T_24; 
  assign _T_72 = _T_71 | _T_32; 
  assign _T_73 = _T_72 | _T_40; 
  assign _T_74 = _T_73 | _T_48; 
  assign _T_75 = _T_74 | _T_56; 
  assign _T_76 = _T_75 | _T_64; 
  assign _T_78 = 23'hff << io_in_a_bits_size; 
  assign _T_79 = _T_78[7:0]; 
  assign _T_80 = ~ _T_79; 
  assign _GEN_33 = {{24'd0}, _T_80}; 
  assign _T_81 = io_in_a_bits_address & _GEN_33; 
  assign _T_82 = _T_81 == 32'h0; 
  assign _T_84 = io_in_a_bits_size[1:0]; 
  assign _T_85 = 4'h1 << _T_84; 
  assign _T_86 = _T_85[2:0]; 
  assign _T_87 = _T_86 | 3'h1; 
  assign _T_88 = io_in_a_bits_size >= 4'h3; 
  assign _T_89 = _T_87[2]; 
  assign _T_90 = io_in_a_bits_address[2]; 
  assign _T_91 = _T_90 == 1'h0; 
  assign _T_93 = _T_89 & _T_91; 
  assign _T_94 = _T_88 | _T_93; 
  assign _T_96 = _T_89 & _T_90; 
  assign _T_97 = _T_88 | _T_96; 
  assign _T_98 = _T_87[1]; 
  assign _T_99 = io_in_a_bits_address[1]; 
  assign _T_100 = _T_99 == 1'h0; 
  assign _T_101 = _T_91 & _T_100; 
  assign _T_102 = _T_98 & _T_101; 
  assign _T_103 = _T_94 | _T_102; 
  assign _T_104 = _T_91 & _T_99; 
  assign _T_105 = _T_98 & _T_104; 
  assign _T_106 = _T_94 | _T_105; 
  assign _T_107 = _T_90 & _T_100; 
  assign _T_108 = _T_98 & _T_107; 
  assign _T_109 = _T_97 | _T_108; 
  assign _T_110 = _T_90 & _T_99; 
  assign _T_111 = _T_98 & _T_110; 
  assign _T_112 = _T_97 | _T_111; 
  assign _T_113 = _T_87[0]; 
  assign _T_114 = io_in_a_bits_address[0]; 
  assign _T_115 = _T_114 == 1'h0; 
  assign _T_116 = _T_101 & _T_115; 
  assign _T_117 = _T_113 & _T_116; 
  assign _T_118 = _T_103 | _T_117; 
  assign _T_119 = _T_101 & _T_114; 
  assign _T_120 = _T_113 & _T_119; 
  assign _T_121 = _T_103 | _T_120; 
  assign _T_122 = _T_104 & _T_115; 
  assign _T_123 = _T_113 & _T_122; 
  assign _T_124 = _T_106 | _T_123; 
  assign _T_125 = _T_104 & _T_114; 
  assign _T_126 = _T_113 & _T_125; 
  assign _T_127 = _T_106 | _T_126; 
  assign _T_128 = _T_107 & _T_115; 
  assign _T_129 = _T_113 & _T_128; 
  assign _T_130 = _T_109 | _T_129; 
  assign _T_131 = _T_107 & _T_114; 
  assign _T_132 = _T_113 & _T_131; 
  assign _T_133 = _T_109 | _T_132; 
  assign _T_134 = _T_110 & _T_115; 
  assign _T_135 = _T_113 & _T_134; 
  assign _T_136 = _T_112 | _T_135; 
  assign _T_137 = _T_110 & _T_114; 
  assign _T_138 = _T_113 & _T_137; 
  assign _T_139 = _T_112 | _T_138; 
  assign _T_146 = {_T_139,_T_136,_T_133,_T_130,_T_127,_T_124,_T_121,_T_118}; 
  assign _T_277 = io_in_a_bits_opcode == 3'h6; 
  assign _T_279 = io_in_a_bits_address ^ 32'h80000000; 
  assign _T_280 = {1'b0,$signed(_T_279)}; 
  assign _T_281 = $signed(_T_280) & $signed(-33'sh80000000); 
  assign _T_282 = $signed(_T_281); 
  assign _T_283 = $signed(_T_282) == $signed(33'sh0); 
  assign _T_284 = io_in_a_bits_address ^ 32'h40000000; 
  assign _T_285 = {1'b0,$signed(_T_284)}; 
  assign _T_286 = $signed(_T_285) & $signed(-33'sh20000000); 
  assign _T_287 = $signed(_T_286); 
  assign _T_288 = $signed(_T_287) == $signed(33'sh0); 
  assign _T_289 = _T_283 | _T_288; 
  assign _T_292 = io_in_a_bits_size <= 4'h6; 
  assign _T_295 = io_in_a_bits_address ^ 32'h10000000; 
  assign _T_296 = {1'b0,$signed(_T_295)}; 
  assign _T_297 = $signed(_T_296) & $signed(-33'sh10000000); 
  assign _T_298 = $signed(_T_297); 
  assign _T_299 = $signed(_T_298) == $signed(33'sh0); 
  assign _T_300 = _T_292 & _T_299; 
  assign _T_304 = _T_300 | reset; 
  assign _T_305 = _T_304 == 1'h0; 
  assign _T_374 = _T_8 ? _T_292 : 1'h0; 
  assign _T_391 = _T_374 | reset; 
  assign _T_392 = _T_391 == 1'h0; 
  assign _T_394 = _T_76 | reset; 
  assign _T_395 = _T_394 == 1'h0; 
  assign _T_398 = _T_88 | reset; 
  assign _T_399 = _T_398 == 1'h0; 
  assign _T_401 = _T_82 | reset; 
  assign _T_402 = _T_401 == 1'h0; 
  assign _T_403 = io_in_a_bits_param <= 3'h2; 
  assign _T_405 = _T_403 | reset; 
  assign _T_406 = _T_405 == 1'h0; 
  assign _T_407 = ~ io_in_a_bits_mask; 
  assign _T_408 = _T_407 == 8'h0; 
  assign _T_410 = _T_408 | reset; 
  assign _T_411 = _T_410 == 1'h0; 
  assign _T_416 = io_in_a_bits_opcode == 3'h7; 
  assign _T_546 = io_in_a_bits_param != 3'h0; 
  assign _T_548 = _T_546 | reset; 
  assign _T_549 = _T_548 == 1'h0; 
  assign _T_559 = io_in_a_bits_opcode == 3'h4; 
  assign _T_580 = _T_289 | _T_299; 
  assign _T_581 = _T_292 & _T_580; 
  assign _T_584 = _T_581 | reset; 
  assign _T_585 = _T_584 == 1'h0; 
  assign _T_592 = io_in_a_bits_param == 3'h0; 
  assign _T_594 = _T_592 | reset; 
  assign _T_595 = _T_594 == 1'h0; 
  assign _T_596 = io_in_a_bits_mask == _T_146; 
  assign _T_598 = _T_596 | reset; 
  assign _T_599 = _T_598 == 1'h0; 
  assign _T_604 = io_in_a_bits_opcode == 3'h0; 
  assign _T_619 = _T_283 | _T_299; 
  assign _T_620 = _T_292 & _T_619; 
  assign _T_622 = io_in_a_bits_size <= 4'h8; 
  assign _T_630 = _T_622 & _T_288; 
  assign _T_632 = _T_620 | _T_630; 
  assign _T_634 = _T_632 | reset; 
  assign _T_635 = _T_634 == 1'h0; 
  assign _T_650 = io_in_a_bits_opcode == 3'h1; 
  assign _T_692 = ~ _T_146; 
  assign _T_693 = io_in_a_bits_mask & _T_692; 
  assign _T_694 = _T_693 == 8'h0; 
  assign _T_696 = _T_694 | reset; 
  assign _T_697 = _T_696 == 1'h0; 
  assign _T_698 = io_in_a_bits_opcode == 3'h2; 
  assign _T_700 = io_in_a_bits_size <= 4'h3; 
  assign _T_720 = _T_700 & _T_580; 
  assign _T_723 = _T_720 | reset; 
  assign _T_724 = _T_723 == 1'h0; 
  assign _T_731 = io_in_a_bits_param <= 3'h4; 
  assign _T_733 = _T_731 | reset; 
  assign _T_734 = _T_733 == 1'h0; 
  assign _T_739 = io_in_a_bits_opcode == 3'h3; 
  assign _T_772 = io_in_a_bits_param <= 3'h3; 
  assign _T_774 = _T_772 | reset; 
  assign _T_775 = _T_774 == 1'h0; 
  assign _T_780 = io_in_a_bits_opcode == 3'h5; 
  assign _T_826 = io_in_d_bits_opcode <= 3'h6; 
  assign _T_828 = _T_826 | reset; 
  assign _T_829 = _T_828 == 1'h0; 
  assign _T_832 = io_in_d_bits_source[5:3]; 
  assign _T_833 = _T_832 == 3'h0; 
  assign _T_841 = _T_832 == 3'h1; 
  assign _T_849 = _T_832 == 3'h2; 
  assign _T_857 = _T_832 == 3'h3; 
  assign _T_865 = _T_832 == 3'h4; 
  assign _T_873 = _T_832 == 3'h5; 
  assign _T_881 = _T_832 == 3'h6; 
  assign _T_889 = _T_832 == 3'h7; 
  assign _T_895 = _T_833 | _T_841; 
  assign _T_896 = _T_895 | _T_849; 
  assign _T_897 = _T_896 | _T_857; 
  assign _T_898 = _T_897 | _T_865; 
  assign _T_899 = _T_898 | _T_873; 
  assign _T_900 = _T_899 | _T_881; 
  assign _T_901 = _T_900 | _T_889; 
  assign _T_902 = io_in_d_bits_sink < 1'h1; 
  assign _T_903 = io_in_d_bits_opcode == 3'h6; 
  assign _T_905 = _T_901 | reset; 
  assign _T_906 = _T_905 == 1'h0; 
  assign _T_907 = io_in_d_bits_size >= 4'h3; 
  assign _T_909 = _T_907 | reset; 
  assign _T_910 = _T_909 == 1'h0; 
  assign _T_911 = io_in_d_bits_param == 2'h0; 
  assign _T_913 = _T_911 | reset; 
  assign _T_914 = _T_913 == 1'h0; 
  assign _T_915 = io_in_d_bits_corrupt == 1'h0; 
  assign _T_917 = _T_915 | reset; 
  assign _T_918 = _T_917 == 1'h0; 
  assign _T_919 = io_in_d_bits_denied == 1'h0; 
  assign _T_921 = _T_919 | reset; 
  assign _T_922 = _T_921 == 1'h0; 
  assign _T_923 = io_in_d_bits_opcode == 3'h4; 
  assign _T_928 = _T_902 | reset; 
  assign _T_929 = _T_928 == 1'h0; 
  assign _T_934 = io_in_d_bits_param <= 2'h2; 
  assign _T_936 = _T_934 | reset; 
  assign _T_937 = _T_936 == 1'h0; 
  assign _T_938 = io_in_d_bits_param != 2'h2; 
  assign _T_940 = _T_938 | reset; 
  assign _T_941 = _T_940 == 1'h0; 
  assign _T_951 = io_in_d_bits_opcode == 3'h5; 
  assign _T_971 = _T_919 | io_in_d_bits_corrupt; 
  assign _T_973 = _T_971 | reset; 
  assign _T_974 = _T_973 == 1'h0; 
  assign _T_980 = io_in_d_bits_opcode == 3'h0; 
  assign _T_997 = io_in_d_bits_opcode == 3'h1; 
  assign _T_1015 = io_in_d_bits_opcode == 3'h2; 
  assign _T_1583 = io_in_c_bits_source[5:3]; 
  assign _T_1584 = _T_1583 == 3'h0; 
  assign _T_1592 = _T_1583 == 3'h1; 
  assign _T_1600 = _T_1583 == 3'h2; 
  assign _T_1608 = _T_1583 == 3'h3; 
  assign _T_1616 = _T_1583 == 3'h4; 
  assign _T_1624 = _T_1583 == 3'h5; 
  assign _T_1632 = _T_1583 == 3'h6; 
  assign _T_1640 = _T_1583 == 3'h7; 
  assign _T_1646 = _T_1584 | _T_1592; 
  assign _T_1647 = _T_1646 | _T_1600; 
  assign _T_1648 = _T_1647 | _T_1608; 
  assign _T_1649 = _T_1648 | _T_1616; 
  assign _T_1650 = _T_1649 | _T_1624; 
  assign _T_1651 = _T_1650 | _T_1632; 
  assign _T_1652 = _T_1651 | _T_1640; 
  assign _T_1654 = 23'hff << io_in_c_bits_size; 
  assign _T_1655 = _T_1654[7:0]; 
  assign _T_1656 = ~ _T_1655; 
  assign _GEN_34 = {{24'd0}, _T_1656}; 
  assign _T_1657 = io_in_c_bits_address & _GEN_34; 
  assign _T_1658 = _T_1657 == 32'h0; 
  assign _T_1659 = io_in_c_bits_address ^ 32'h80000000; 
  assign _T_1660 = {1'b0,$signed(_T_1659)}; 
  assign _T_1661 = $signed(_T_1660) & $signed(-33'sh80000000); 
  assign _T_1662 = $signed(_T_1661); 
  assign _T_1663 = $signed(_T_1662) == $signed(33'sh0); 
  assign _T_1664 = io_in_c_bits_address ^ 32'h40000000; 
  assign _T_1665 = {1'b0,$signed(_T_1664)}; 
  assign _T_1666 = $signed(_T_1665) & $signed(-33'sh20000000); 
  assign _T_1667 = $signed(_T_1666); 
  assign _T_1668 = $signed(_T_1667) == $signed(33'sh0); 
  assign _T_1669 = io_in_c_bits_address ^ 32'h10000000; 
  assign _T_1670 = {1'b0,$signed(_T_1669)}; 
  assign _T_1671 = $signed(_T_1670) & $signed(-33'sh10000000); 
  assign _T_1672 = $signed(_T_1671); 
  assign _T_1673 = $signed(_T_1672) == $signed(33'sh0); 
  assign _T_1675 = _T_1663 | _T_1668; 
  assign _T_1676 = _T_1675 | _T_1673; 
  assign _T_1807 = io_in_c_bits_opcode == 3'h4; 
  assign _T_1809 = _T_1676 | reset; 
  assign _T_1810 = _T_1809 == 1'h0; 
  assign _T_1812 = _T_1652 | reset; 
  assign _T_1813 = _T_1812 == 1'h0; 
  assign _T_1814 = io_in_c_bits_size >= 4'h3; 
  assign _T_1816 = _T_1814 | reset; 
  assign _T_1817 = _T_1816 == 1'h0; 
  assign _T_1819 = _T_1658 | reset; 
  assign _T_1820 = _T_1819 == 1'h0; 
  assign _T_1821 = io_in_c_bits_param <= 3'h5; 
  assign _T_1823 = _T_1821 | reset; 
  assign _T_1824 = _T_1823 == 1'h0; 
  assign _T_1825 = io_in_c_bits_corrupt == 1'h0; 
  assign _T_1827 = _T_1825 | reset; 
  assign _T_1828 = _T_1827 == 1'h0; 
  assign _T_1829 = io_in_c_bits_opcode == 3'h5; 
  assign _T_1847 = io_in_c_bits_opcode == 3'h6; 
  assign _T_1862 = io_in_c_bits_size <= 4'h6; 
  assign _T_1870 = _T_1862 & _T_1673; 
  assign _T_1874 = _T_1870 | reset; 
  assign _T_1875 = _T_1874 == 1'h0; 
  assign _T_1944 = _T_1584 ? _T_1862 : 1'h0; 
  assign _T_1961 = _T_1944 | reset; 
  assign _T_1962 = _T_1961 == 1'h0; 
  assign _T_1973 = io_in_c_bits_param <= 3'h2; 
  assign _T_1975 = _T_1973 | reset; 
  assign _T_1976 = _T_1975 == 1'h0; 
  assign _T_1981 = io_in_c_bits_opcode == 3'h7; 
  assign _T_2111 = io_in_c_bits_opcode == 3'h0; 
  assign _T_2121 = io_in_c_bits_param == 3'h0; 
  assign _T_2123 = _T_2121 | reset; 
  assign _T_2124 = _T_2123 == 1'h0; 
  assign _T_2129 = io_in_c_bits_opcode == 3'h1; 
  assign _T_2143 = io_in_c_bits_opcode == 3'h2; 
  assign _T_2161 = io_in_e_bits_sink < 1'h1; 
  assign _T_2163 = _T_2161 | reset; 
  assign _T_2164 = _T_2163 == 1'h0; 
  assign _T_2165 = io_in_a_ready & io_in_a_valid; 
  assign _T_2170 = _T_80[7:3]; 
  assign _T_2171 = io_in_a_bits_opcode[2]; 
  assign _T_2172 = _T_2171 == 1'h0; 
  assign _T_2176 = _T_2174 - 5'h1; 
  assign _T_2177 = _T_2174 == 5'h0; 
  assign _T_2190 = _T_2177 == 1'h0; 
  assign _T_2191 = io_in_a_valid & _T_2190; 
  assign _T_2192 = io_in_a_bits_opcode == _T_2185; 
  assign _T_2194 = _T_2192 | reset; 
  assign _T_2195 = _T_2194 == 1'h0; 
  assign _T_2196 = io_in_a_bits_param == _T_2186; 
  assign _T_2198 = _T_2196 | reset; 
  assign _T_2199 = _T_2198 == 1'h0; 
  assign _T_2200 = io_in_a_bits_size == _T_2187; 
  assign _T_2202 = _T_2200 | reset; 
  assign _T_2203 = _T_2202 == 1'h0; 
  assign _T_2204 = io_in_a_bits_source == _T_2188; 
  assign _T_2206 = _T_2204 | reset; 
  assign _T_2207 = _T_2206 == 1'h0; 
  assign _T_2208 = io_in_a_bits_address == _T_2189; 
  assign _T_2210 = _T_2208 | reset; 
  assign _T_2211 = _T_2210 == 1'h0; 
  assign _T_2213 = _T_2165 & _T_2177; 
  assign _T_2214 = io_in_d_ready & io_in_d_valid; 
  assign _T_2216 = 23'hff << io_in_d_bits_size; 
  assign _T_2217 = _T_2216[7:0]; 
  assign _T_2218 = ~ _T_2217; 
  assign _T_2219 = _T_2218[7:3]; 
  assign _T_2220 = io_in_d_bits_opcode[0]; 
  assign _T_2224 = _T_2222 - 5'h1; 
  assign _T_2225 = _T_2222 == 5'h0; 
  assign _T_2239 = _T_2225 == 1'h0; 
  assign _T_2240 = io_in_d_valid & _T_2239; 
  assign _T_2241 = io_in_d_bits_opcode == _T_2233; 
  assign _T_2243 = _T_2241 | reset; 
  assign _T_2244 = _T_2243 == 1'h0; 
  assign _T_2245 = io_in_d_bits_param == _T_2234; 
  assign _T_2247 = _T_2245 | reset; 
  assign _T_2248 = _T_2247 == 1'h0; 
  assign _T_2249 = io_in_d_bits_size == _T_2235; 
  assign _T_2251 = _T_2249 | reset; 
  assign _T_2252 = _T_2251 == 1'h0; 
  assign _T_2253 = io_in_d_bits_source == _T_2236; 
  assign _T_2255 = _T_2253 | reset; 
  assign _T_2256 = _T_2255 == 1'h0; 
  assign _T_2257 = io_in_d_bits_sink == _T_2237; 
  assign _T_2259 = _T_2257 | reset; 
  assign _T_2260 = _T_2259 == 1'h0; 
  assign _T_2261 = io_in_d_bits_denied == _T_2238; 
  assign _T_2263 = _T_2261 | reset; 
  assign _T_2264 = _T_2263 == 1'h0; 
  assign _T_2266 = _T_2214 & _T_2225; 
  assign _T_2316 = io_in_c_ready & io_in_c_valid; 
  assign _T_2321 = _T_1656[7:3]; 
  assign _T_2322 = io_in_c_bits_opcode[0]; 
  assign _T_2326 = _T_2324 - 5'h1; 
  assign _T_2327 = _T_2324 == 5'h0; 
  assign _T_2340 = _T_2327 == 1'h0; 
  assign _T_2341 = io_in_c_valid & _T_2340; 
  assign _T_2342 = io_in_c_bits_opcode == _T_2335; 
  assign _T_2344 = _T_2342 | reset; 
  assign _T_2345 = _T_2344 == 1'h0; 
  assign _T_2346 = io_in_c_bits_param == _T_2336; 
  assign _T_2348 = _T_2346 | reset; 
  assign _T_2349 = _T_2348 == 1'h0; 
  assign _T_2350 = io_in_c_bits_size == _T_2337; 
  assign _T_2352 = _T_2350 | reset; 
  assign _T_2353 = _T_2352 == 1'h0; 
  assign _T_2354 = io_in_c_bits_source == _T_2338; 
  assign _T_2356 = _T_2354 | reset; 
  assign _T_2357 = _T_2356 == 1'h0; 
  assign _T_2358 = io_in_c_bits_address == _T_2339; 
  assign _T_2360 = _T_2358 | reset; 
  assign _T_2361 = _T_2360 == 1'h0; 
  assign _T_2363 = _T_2316 & _T_2327; 
  assign _T_2376 = _T_2374 - 5'h1; 
  assign _T_2377 = _T_2374 == 5'h0; 
  assign _T_2395 = _T_2393 - 5'h1; 
  assign _T_2396 = _T_2393 == 5'h0; 
  assign _T_2406 = _T_2165 & _T_2377; 
  assign _T_2408 = 64'h1 << io_in_a_bits_source; 
  assign _T_2409 = _T_2364 >> io_in_a_bits_source; 
  assign _T_2410 = _T_2409[0]; 
  assign _T_2411 = _T_2410 == 1'h0; 
  assign _T_2413 = _T_2411 | reset; 
  assign _T_2414 = _T_2413 == 1'h0; 
  assign _GEN_27 = _T_2406 ? _T_2408 : 64'h0; 
  assign _T_2418 = _T_2214 & _T_2396; 
  assign _T_2420 = _T_903 == 1'h0; 
  assign _T_2421 = _T_2418 & _T_2420; 
  assign _T_2422 = 64'h1 << io_in_d_bits_source; 
  assign _T_2423 = _GEN_27 | _T_2364; 
  assign _T_2424 = _T_2423 >> io_in_d_bits_source; 
  assign _T_2425 = _T_2424[0]; 
  assign _T_2427 = _T_2425 | reset; 
  assign _T_2428 = _T_2427 == 1'h0; 
  assign _GEN_28 = _T_2421 ? _T_2422 : 64'h0; 
  assign _T_2429 = _GEN_27 != _GEN_28; 
  assign _T_2430 = _GEN_27 != 64'h0; 
  assign _T_2431 = _T_2430 == 1'h0; 
  assign _T_2432 = _T_2429 | _T_2431; 
  assign _T_2434 = _T_2432 | reset; 
  assign _T_2435 = _T_2434 == 1'h0; 
  assign _T_2436 = _T_2364 | _GEN_27; 
  assign _T_2437 = ~ _GEN_28; 
  assign _T_2438 = _T_2436 & _T_2437; 
  assign _T_2440 = _T_2364 != 64'h0; 
  assign _T_2441 = _T_2440 == 1'h0; 
  assign _T_2442 = plusarg_reader_out == 32'h0; 
  assign _T_2443 = _T_2441 | _T_2442; 
  assign _T_2444 = _T_2439 < plusarg_reader_out; 
  assign _T_2445 = _T_2443 | _T_2444; 
  assign _T_2447 = _T_2445 | reset; 
  assign _T_2448 = _T_2447 == 1'h0; 
  assign _T_2450 = _T_2439 + 32'h1; 
  assign _T_2453 = _T_2165 | _T_2214; 
  assign _T_2465 = _T_2463 - 5'h1; 
  assign _T_2466 = _T_2463 == 5'h0; 
  assign _T_2476 = _T_2214 & _T_2466; 
  assign _T_2477 = io_in_d_bits_opcode[2]; 
  assign _T_2478 = io_in_d_bits_opcode[1]; 
  assign _T_2479 = _T_2478 == 1'h0; 
  assign _T_2480 = _T_2477 & _T_2479; 
  assign _T_2481 = _T_2476 & _T_2480; 
  assign _T_2482 = 2'h1 << io_in_d_bits_sink; 
  assign _T_2483 = _T_2454 >> io_in_d_bits_sink; 
  assign _T_2485 = _T_2483 == 1'h0; 
  assign _T_2487 = _T_2485 | reset; 
  assign _T_2488 = _T_2487 == 1'h0; 
  assign _GEN_31 = _T_2481 ? _T_2482 : 2'h0; 
  assign _T_2490 = io_in_e_ready & io_in_e_valid; 
  assign _T_2493 = 2'h1 << io_in_e_bits_sink; 
  assign _T_2474 = _GEN_31[0]; 
  assign _T_2494 = _T_2474 | _T_2454; 
  assign _T_2495 = _T_2494 >> io_in_e_bits_sink; 
  assign _T_2498 = _T_2495 | reset; 
  assign _T_2499 = _T_2498 == 1'h0; 
  assign _GEN_32 = _T_2490 ? _T_2493 : 2'h0; 
  assign _T_2500 = _T_2454 | _T_2474; 
  assign _T_2489 = _GEN_32[0]; 
  assign _T_2501 = ~ _T_2489; 
  assign _T_2502 = _T_2500 & _T_2501; 
  assign _GEN_35 = io_in_a_valid & _T_277; 
  assign _GEN_49 = io_in_a_valid & _T_416; 
  assign _GEN_65 = io_in_a_valid & _T_559; 
  assign _GEN_75 = io_in_a_valid & _T_604; 
  assign _GEN_85 = io_in_a_valid & _T_650; 
  assign _GEN_95 = io_in_a_valid & _T_698; 
  assign _GEN_105 = io_in_a_valid & _T_739; 
  assign _GEN_115 = io_in_a_valid & _T_780; 
  assign _GEN_123 = io_in_d_valid & _T_903; 
  assign _GEN_133 = io_in_d_valid & _T_923; 
  assign _GEN_145 = io_in_d_valid & _T_951; 
  assign _GEN_157 = io_in_d_valid & _T_980; 
  assign _GEN_163 = io_in_d_valid & _T_997; 
  assign _GEN_169 = io_in_d_valid & _T_1015; 
  assign _GEN_175 = io_in_c_valid & _T_1807; 
  assign _GEN_187 = io_in_c_valid & _T_1829; 
  assign _GEN_197 = io_in_c_valid & _T_1847; 
  assign _GEN_211 = io_in_c_valid & _T_1981; 
  assign _GEN_223 = io_in_c_valid & _T_2111; 
  assign _GEN_233 = io_in_c_valid & _T_2129; 
  assign _GEN_241 = io_in_c_valid & _T_2143; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2174 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_2185 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2186 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_2187 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_2188 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_2189 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_2222 = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_2233 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_2234 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_2235 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_2236 = _RAND_10[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_2237 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_2238 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_2324 = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_2335 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_2336 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_2337 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_2338 = _RAND_17[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_2339 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  _T_2364 = _RAND_19[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_2374 = _RAND_20[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_2393 = _RAND_21[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_2439 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_2454 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_2463 = _RAND_24[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_2174 <= 5'h0;
    end else begin
      if (_T_2165) begin
        if (_T_2177) begin
          if (_T_2172) begin
            _T_2174 <= _T_2170;
          end else begin
            _T_2174 <= 5'h0;
          end
        end else begin
          _T_2174 <= _T_2176;
        end
      end
    end
    if (_T_2213) begin
      _T_2185 <= io_in_a_bits_opcode;
    end
    if (_T_2213) begin
      _T_2186 <= io_in_a_bits_param;
    end
    if (_T_2213) begin
      _T_2187 <= io_in_a_bits_size;
    end
    if (_T_2213) begin
      _T_2188 <= io_in_a_bits_source;
    end
    if (_T_2213) begin
      _T_2189 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_2222 <= 5'h0;
    end else begin
      if (_T_2214) begin
        if (_T_2225) begin
          if (_T_2220) begin
            _T_2222 <= _T_2219;
          end else begin
            _T_2222 <= 5'h0;
          end
        end else begin
          _T_2222 <= _T_2224;
        end
      end
    end
    if (_T_2266) begin
      _T_2233 <= io_in_d_bits_opcode;
    end
    if (_T_2266) begin
      _T_2234 <= io_in_d_bits_param;
    end
    if (_T_2266) begin
      _T_2235 <= io_in_d_bits_size;
    end
    if (_T_2266) begin
      _T_2236 <= io_in_d_bits_source;
    end
    if (_T_2266) begin
      _T_2237 <= io_in_d_bits_sink;
    end
    if (_T_2266) begin
      _T_2238 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_2324 <= 5'h0;
    end else begin
      if (_T_2316) begin
        if (_T_2327) begin
          if (_T_2322) begin
            _T_2324 <= _T_2321;
          end else begin
            _T_2324 <= 5'h0;
          end
        end else begin
          _T_2324 <= _T_2326;
        end
      end
    end
    if (_T_2363) begin
      _T_2335 <= io_in_c_bits_opcode;
    end
    if (_T_2363) begin
      _T_2336 <= io_in_c_bits_param;
    end
    if (_T_2363) begin
      _T_2337 <= io_in_c_bits_size;
    end
    if (_T_2363) begin
      _T_2338 <= io_in_c_bits_source;
    end
    if (_T_2363) begin
      _T_2339 <= io_in_c_bits_address;
    end
    if (reset) begin
      _T_2364 <= 64'h0;
    end else begin
      _T_2364 <= _T_2438;
    end
    if (reset) begin
      _T_2374 <= 5'h0;
    end else begin
      if (_T_2165) begin
        if (_T_2377) begin
          if (_T_2172) begin
            _T_2374 <= _T_2170;
          end else begin
            _T_2374 <= 5'h0;
          end
        end else begin
          _T_2374 <= _T_2376;
        end
      end
    end
    if (reset) begin
      _T_2393 <= 5'h0;
    end else begin
      if (_T_2214) begin
        if (_T_2396) begin
          if (_T_2220) begin
            _T_2393 <= _T_2219;
          end else begin
            _T_2393 <= 5'h0;
          end
        end else begin
          _T_2393 <= _T_2395;
        end
      end
    end
    if (reset) begin
      _T_2439 <= 32'h0;
    end else begin
      if (_T_2453) begin
        _T_2439 <= 32'h0;
      end else begin
        _T_2439 <= _T_2450;
      end
    end
    if (reset) begin
      _T_2454 <= 1'h0;
    end else begin
      _T_2454 <= _T_2502;
    end
    if (reset) begin
      _T_2463 <= 5'h0;
    end else begin
      if (_T_2214) begin
        if (_T_2466) begin
          if (_T_2220) begin
            _T_2463 <= _T_2219;
          end else begin
            _T_2463 <= 5'h0;
          end
        end else begin
          _T_2463 <= _T_2465;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel has invalid opcode (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:39 assert (TLMessages.isA(bundle.opcode), \"'A' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:46 assert (visible(edge.address(bundle), bundle.source, edge), \"'A' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_305) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_305) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_392) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_392) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_399) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_399) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_406) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_406) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_411) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_411) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:56 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_305) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_305) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_392) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_392) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_399) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_399) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_406) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_406) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_549) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_549) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_411) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_411) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:68 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_585) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_585) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_595) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_595) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_599) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:77 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_635) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_635) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_595) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_595) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_599) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_635) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_635) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_595) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_595) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_697) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_697) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_724) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_724) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_734) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_734) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_599) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_724) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_724) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_775) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_775) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_599) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_635) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_635) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_599) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:117 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_829) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_829) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_906) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_906) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_910) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_910) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_914) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_914) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_918) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_918) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_922) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_922) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_906) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_906) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_929) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:285 assert (sink_ok, \"'D' channel Grant carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_929) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_910) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_910) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_937) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_937) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_941) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_941) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_918) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_918) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is denied (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:290 assert (deny_put_ok || !bundle.denied, \"'D' channel Grant is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_906) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_906) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_929) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:295 assert (sink_ok, \"'D' channel GrantData carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_929) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_910) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_910) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_937) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_937) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_941) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_941) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_974) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_974) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:300 assert (deny_get_ok || !bundle.denied, \"'D' channel GrantData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_157 & _T_906) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_157 & _T_906) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_157 & _T_914) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_157 & _T_914) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_157 & _T_918) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_157 & _T_918) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is denied (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:308 assert (deny_put_ok || !bundle.denied, \"'D' channel AccessAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_906) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_906) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_914) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_914) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_974) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_974) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:316 assert (deny_get_ok || !bundle.denied, \"'D' channel AccessAckData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_169 & _T_906) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_169 & _T_906) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_169 & _T_914) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_169 & _T_914) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_169 & _T_918) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_169 & _T_918) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is denied (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:324 assert (deny_put_ok || !bundle.denied, \"'D' channel HintAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel has invalid opcode (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:122 assert (TLMessages.isB(bundle.opcode), \"'B' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:124 assert (visible(edge.address(bundle), bundle.source, edge), \"'B' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Probe type unsupported by client (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:133 assert (edge.client.supportsProbe(bundle.source, bundle.size), \"'B' channel carries Probe type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:134 assert (address_ok, \"'B' channel Probe carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries source that is not first source (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:135 assert (legal_source, \"'B' channel Probe carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:136 assert (is_aligned, \"'B' channel Probe address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:137 assert (TLPermissions.isCap(bundle.param), \"'B' channel Probe carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe contains invalid mask (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:138 assert (bundle.mask === mask, \"'B' channel Probe contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe is corrupt (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:139 assert (!bundle.corrupt, \"'B' channel Probe is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Get type unsupported by client (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:143 assert (edge.client.supportsGet(bundle.source, bundle.size), \"'B' channel carries Get type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries unmanaged address (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:144 assert (address_ok, \"'B' channel Get carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries source that is not first source (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:145 assert (legal_source, \"'B' channel Get carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:146 assert (is_aligned, \"'B' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries invalid param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:147 assert (bundle.param === UInt(0), \"'B' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get contains invalid mask (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:148 assert (bundle.mask === mask, \"'B' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get is corrupt (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:149 assert (!bundle.corrupt, \"'B' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutFull type unsupported by client (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:153 assert (edge.client.supportsPutFull(bundle.source, bundle.size), \"'B' channel carries PutFull type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries unmanaged address (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:154 assert (address_ok, \"'B' channel PutFull carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries source that is not first source (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:155 assert (legal_source, \"'B' channel PutFull carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:156 assert (is_aligned, \"'B' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries invalid param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:157 assert (bundle.param === UInt(0), \"'B' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull contains invalid mask (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:158 assert (bundle.mask === mask, \"'B' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutPartial type unsupported by client (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:162 assert (edge.client.supportsPutPartial(bundle.source, bundle.size), \"'B' channel carries PutPartial type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:163 assert (address_ok, \"'B' channel PutPartial carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:164 assert (legal_source, \"'B' channel PutPartial carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:165 assert (is_aligned, \"'B' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries invalid param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:166 assert (bundle.param === UInt(0), \"'B' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial contains invalid mask (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:167 assert ((bundle.mask & ~mask) === UInt(0), \"'B' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Arithmetic type unsupported by client (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:171 assert (edge.client.supportsArithmetic(bundle.source, bundle.size), \"'B' channel carries Arithmetic type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:172 assert (address_ok, \"'B' channel Arithmetic carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:173 assert (legal_source, \"'B' channel Arithmetic carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:174 assert (is_aligned, \"'B' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries invalid opcode param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:175 assert (TLAtomics.isArithmetic(bundle.param), \"'B' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:176 assert (bundle.mask === mask, \"'B' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Logical type unsupported by client (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:180 assert (edge.client.supportsLogical(bundle.source, bundle.size), \"'B' channel carries Logical type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries unmanaged address (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:181 assert (address_ok, \"'B' channel Logical carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries source that is not first source (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:182 assert (legal_source, \"'B' channel Logical carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:183 assert (is_aligned, \"'B' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries invalid opcode param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:184 assert (TLAtomics.isLogical(bundle.param), \"'B' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical contains invalid mask (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:185 assert (bundle.mask === mask, \"'B' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Hint type unsupported by client (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:189 assert (edge.client.supportsHint(bundle.source, bundle.size), \"'B' channel carries Hint type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries unmanaged address (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:190 assert (address_ok, \"'B' channel Hint carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries source that is not first source (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:191 assert (legal_source, \"'B' channel Hint carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:192 assert (is_aligned, \"'B' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint contains invalid mask (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:193 assert (bundle.mask === mask, \"'B' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint is corrupt (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:194 assert (!bundle.corrupt, \"'B' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel has invalid opcode (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:199 assert (TLMessages.isC(bundle.opcode), \"'C' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:205 assert (visible(edge.address(bundle), bundle.source, edge), \"'C' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1810) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:208 assert (address_ok, \"'C' channel ProbeAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1810) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1813) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:209 assert (source_ok, \"'C' channel ProbeAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1813) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1817) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:210 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1817) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1820) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:211 assert (is_aligned, \"'C' channel ProbeAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1820) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1824) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:212 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAck carries invalid report param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1824) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1828) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck is corrupt (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:213 assert (!bundle.corrupt, \"'C' channel ProbeAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1828) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_187 & _T_1810) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:217 assert (address_ok, \"'C' channel ProbeAckData carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_187 & _T_1810) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_187 & _T_1813) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:218 assert (source_ok, \"'C' channel ProbeAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_187 & _T_1813) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_187 & _T_1817) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:219 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAckData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_187 & _T_1817) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_187 & _T_1820) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:220 assert (is_aligned, \"'C' channel ProbeAckData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_187 & _T_1820) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_187 & _T_1824) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:221 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAckData carries invalid report param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_187 & _T_1824) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1875) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:225 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries Release type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1875) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1962) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:226 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1962) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1813) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:227 assert (source_ok, \"'C' channel Release carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1813) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1817) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:228 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel Release smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1817) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1820) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:229 assert (is_aligned, \"'C' channel Release address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1820) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1976) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid shrink param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:230 assert (TLPermissions.isShrink(bundle.param), \"'C' channel Release carries invalid shrink param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1976) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1828) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release is corrupt (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:231 assert (!bundle.corrupt, \"'C' channel Release is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1828) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1875) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:235 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries ReleaseData type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1875) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1962) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:236 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1962) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1813) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:237 assert (source_ok, \"'C' channel ReleaseData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1813) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1817) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:238 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ReleaseData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1817) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1820) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:239 assert (is_aligned, \"'C' channel ReleaseData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1820) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1976) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid shrink param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:240 assert (TLPermissions.isShrink(bundle.param), \"'C' channel ReleaseData carries invalid shrink param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1976) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_1810) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:244 assert (address_ok, \"'C' channel AccessAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_1810) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_1813) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:245 assert (source_ok, \"'C' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_1813) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_1820) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:246 assert (is_aligned, \"'C' channel AccessAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_1820) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_2124) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:247 assert (bundle.param === UInt(0), \"'C' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_2124) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_1828) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck is corrupt (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:248 assert (!bundle.corrupt, \"'C' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_1828) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_1810) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:252 assert (address_ok, \"'C' channel AccessAckData carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_1810) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_1813) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:253 assert (source_ok, \"'C' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_1813) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_1820) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:254 assert (is_aligned, \"'C' channel AccessAckData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_1820) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_2124) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:255 assert (bundle.param === UInt(0), \"'C' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_2124) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1810) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:259 assert (address_ok, \"'C' channel HintAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1810) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1813) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:260 assert (source_ok, \"'C' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1813) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1820) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:261 assert (is_aligned, \"'C' channel HintAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1820) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_2124) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:262 assert (bundle.param === UInt(0), \"'C' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_2124) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1828) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck is corrupt (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:263 assert (!bundle.corrupt, \"'C' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1828) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_e_valid & _T_2164) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channels carries invalid sink ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:330 assert (sink_ok, \"'E' channels carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_e_valid & _T_2164) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2191 & _T_2195) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2191 & _T_2195) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2191 & _T_2199) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2191 & _T_2199) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2191 & _T_2203) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2191 & _T_2203) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2191 & _T_2207) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2191 & _T_2207) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2191 & _T_2211) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2191 & _T_2211) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2240 & _T_2244) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2240 & _T_2244) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2240 & _T_2248) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2240 & _T_2248) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2240 & _T_2252) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2240 & _T_2252) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2240 & _T_2256) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2240 & _T_2256) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2240 & _T_2260) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2240 & _T_2260) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2240 & _T_2264) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2240 & _T_2264) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:378 assert (b.bits.opcode === opcode, \"'B' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:379 assert (b.bits.param  === param,  \"'B' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel size changed within multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:380 assert (b.bits.size   === size,   \"'B' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel source changed within multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:381 assert (b.bits.source === source, \"'B' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:382 assert (b.bits.address=== address,\"'B' channel addresss changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2341 & _T_2345) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:401 assert (c.bits.opcode === opcode, \"'C' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2341 & _T_2345) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2341 & _T_2349) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:402 assert (c.bits.param  === param,  \"'C' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2341 & _T_2349) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2341 & _T_2353) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:403 assert (c.bits.size   === size,   \"'C' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2341 & _T_2353) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2341 & _T_2357) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:404 assert (c.bits.source === source, \"'C' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2341 & _T_2357) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2341 & _T_2361) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:405 assert (c.bits.address=== address,\"'C' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2341 & _T_2361) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2406 & _T_2414) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2406 & _T_2414) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2421 & _T_2428) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2421 & _T_2428) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2435) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2435) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2448) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:479 assert (!inflight.orR || limit === UInt(0) || watchdog < limit, \"TileLink timeout expired\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2448) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2481 & _T_2488) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:494 assert(!inflight(bundle.d.bits.sink), \"'D' channel re-used a sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2481 & _T_2488) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2490 & _T_2499) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at ChiplinkTest.scala:362:98)\n    at Monitor.scala:500 assert((d_set | inflight)(bundle.e.bits.sink), \"'E' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2490 & _T_2499) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLMonitor_17( 
  input         clock, 
  input         reset, 
  input         io_in_a_ready, 
  input         io_in_a_valid, 
  input  [2:0]  io_in_a_bits_opcode, 
  input  [2:0]  io_in_a_bits_param, 
  input  [3:0]  io_in_a_bits_size, 
  input  [5:0]  io_in_a_bits_source, 
  input  [31:0] io_in_a_bits_address, 
  input  [3:0]  io_in_a_bits_mask, 
  input         io_in_c_ready, 
  input         io_in_c_valid, 
  input  [2:0]  io_in_c_bits_opcode, 
  input  [2:0]  io_in_c_bits_param, 
  input  [3:0]  io_in_c_bits_size, 
  input  [5:0]  io_in_c_bits_source, 
  input  [31:0] io_in_c_bits_address, 
  input         io_in_c_bits_corrupt, 
  input         io_in_d_ready, 
  input         io_in_d_valid, 
  input  [2:0]  io_in_d_bits_opcode, 
  input  [1:0]  io_in_d_bits_param, 
  input  [3:0]  io_in_d_bits_size, 
  input  [5:0]  io_in_d_bits_source, 
  input         io_in_d_bits_sink, 
  input         io_in_d_bits_denied, 
  input         io_in_d_bits_corrupt, 
  input         io_in_e_ready, 
  input         io_in_e_valid, 
  input         io_in_e_bits_sink 
);
  wire [31:0] plusarg_reader_out; 
  wire [2:0] _T_7; 
  wire  _T_8; 
  wire  _T_16; 
  wire  _T_24; 
  wire  _T_32; 
  wire  _T_40; 
  wire  _T_48; 
  wire  _T_56; 
  wire  _T_64; 
  wire  _T_70; 
  wire  _T_71; 
  wire  _T_72; 
  wire  _T_73; 
  wire  _T_74; 
  wire  _T_75; 
  wire  _T_76; 
  wire [22:0] _T_78; 
  wire [7:0] _T_79; 
  wire [7:0] _T_80; 
  wire [31:0] _GEN_33; 
  wire [31:0] _T_81; 
  wire  _T_82; 
  wire  _T_84; 
  wire [1:0] _T_85; 
  wire [1:0] _T_87; 
  wire  _T_88; 
  wire  _T_89; 
  wire  _T_90; 
  wire  _T_91; 
  wire  _T_93; 
  wire  _T_94; 
  wire  _T_96; 
  wire  _T_97; 
  wire  _T_98; 
  wire  _T_99; 
  wire  _T_100; 
  wire  _T_101; 
  wire  _T_102; 
  wire  _T_103; 
  wire  _T_104; 
  wire  _T_105; 
  wire  _T_106; 
  wire  _T_107; 
  wire  _T_108; 
  wire  _T_109; 
  wire  _T_110; 
  wire  _T_111; 
  wire  _T_112; 
  wire [3:0] _T_115; 
  wire  _T_246; 
  wire [31:0] _T_248; 
  wire [32:0] _T_249; 
  wire [32:0] _T_250; 
  wire [32:0] _T_251; 
  wire  _T_252; 
  wire [31:0] _T_253; 
  wire [32:0] _T_254; 
  wire [32:0] _T_255; 
  wire [32:0] _T_256; 
  wire  _T_257; 
  wire  _T_258; 
  wire  _T_261; 
  wire [31:0] _T_264; 
  wire [32:0] _T_265; 
  wire [32:0] _T_266; 
  wire [32:0] _T_267; 
  wire  _T_268; 
  wire  _T_269; 
  wire  _T_273; 
  wire  _T_274; 
  wire  _T_343; 
  wire  _T_360; 
  wire  _T_361; 
  wire  _T_363; 
  wire  _T_364; 
  wire  _T_367; 
  wire  _T_368; 
  wire  _T_370; 
  wire  _T_371; 
  wire  _T_372; 
  wire  _T_374; 
  wire  _T_375; 
  wire [3:0] _T_376; 
  wire  _T_377; 
  wire  _T_379; 
  wire  _T_380; 
  wire  _T_385; 
  wire  _T_515; 
  wire  _T_517; 
  wire  _T_518; 
  wire  _T_528; 
  wire  _T_549; 
  wire  _T_550; 
  wire  _T_553; 
  wire  _T_554; 
  wire  _T_561; 
  wire  _T_563; 
  wire  _T_564; 
  wire  _T_565; 
  wire  _T_567; 
  wire  _T_568; 
  wire  _T_573; 
  wire  _T_588; 
  wire  _T_589; 
  wire  _T_591; 
  wire  _T_599; 
  wire  _T_601; 
  wire  _T_603; 
  wire  _T_604; 
  wire  _T_619; 
  wire [3:0] _T_661; 
  wire [3:0] _T_662; 
  wire  _T_663; 
  wire  _T_665; 
  wire  _T_666; 
  wire  _T_667; 
  wire  _T_669; 
  wire  _T_689; 
  wire  _T_692; 
  wire  _T_693; 
  wire  _T_700; 
  wire  _T_702; 
  wire  _T_703; 
  wire  _T_708; 
  wire  _T_741; 
  wire  _T_743; 
  wire  _T_744; 
  wire  _T_749; 
  wire  _T_795; 
  wire  _T_797; 
  wire  _T_798; 
  wire [2:0] _T_801; 
  wire  _T_802; 
  wire  _T_810; 
  wire  _T_818; 
  wire  _T_826; 
  wire  _T_834; 
  wire  _T_842; 
  wire  _T_850; 
  wire  _T_858; 
  wire  _T_864; 
  wire  _T_865; 
  wire  _T_866; 
  wire  _T_867; 
  wire  _T_868; 
  wire  _T_869; 
  wire  _T_870; 
  wire  _T_871; 
  wire  _T_872; 
  wire  _T_874; 
  wire  _T_875; 
  wire  _T_876; 
  wire  _T_878; 
  wire  _T_879; 
  wire  _T_880; 
  wire  _T_882; 
  wire  _T_883; 
  wire  _T_884; 
  wire  _T_886; 
  wire  _T_887; 
  wire  _T_888; 
  wire  _T_890; 
  wire  _T_891; 
  wire  _T_892; 
  wire  _T_897; 
  wire  _T_898; 
  wire  _T_903; 
  wire  _T_905; 
  wire  _T_906; 
  wire  _T_907; 
  wire  _T_909; 
  wire  _T_910; 
  wire  _T_920; 
  wire  _T_940; 
  wire  _T_942; 
  wire  _T_943; 
  wire  _T_949; 
  wire  _T_966; 
  wire  _T_984; 
  wire [2:0] _T_1521; 
  wire  _T_1522; 
  wire  _T_1530; 
  wire  _T_1538; 
  wire  _T_1546; 
  wire  _T_1554; 
  wire  _T_1562; 
  wire  _T_1570; 
  wire  _T_1578; 
  wire  _T_1584; 
  wire  _T_1585; 
  wire  _T_1586; 
  wire  _T_1587; 
  wire  _T_1588; 
  wire  _T_1589; 
  wire  _T_1590; 
  wire [22:0] _T_1592; 
  wire [7:0] _T_1593; 
  wire [7:0] _T_1594; 
  wire [31:0] _GEN_34; 
  wire [31:0] _T_1595; 
  wire  _T_1596; 
  wire [31:0] _T_1597; 
  wire [32:0] _T_1598; 
  wire [32:0] _T_1599; 
  wire [32:0] _T_1600; 
  wire  _T_1601; 
  wire [31:0] _T_1602; 
  wire [32:0] _T_1603; 
  wire [32:0] _T_1604; 
  wire [32:0] _T_1605; 
  wire  _T_1606; 
  wire [31:0] _T_1607; 
  wire [32:0] _T_1608; 
  wire [32:0] _T_1609; 
  wire [32:0] _T_1610; 
  wire  _T_1611; 
  wire  _T_1613; 
  wire  _T_1614; 
  wire  _T_1745; 
  wire  _T_1747; 
  wire  _T_1748; 
  wire  _T_1750; 
  wire  _T_1751; 
  wire  _T_1752; 
  wire  _T_1754; 
  wire  _T_1755; 
  wire  _T_1757; 
  wire  _T_1758; 
  wire  _T_1759; 
  wire  _T_1761; 
  wire  _T_1762; 
  wire  _T_1763; 
  wire  _T_1765; 
  wire  _T_1766; 
  wire  _T_1767; 
  wire  _T_1785; 
  wire  _T_1800; 
  wire  _T_1808; 
  wire  _T_1812; 
  wire  _T_1813; 
  wire  _T_1882; 
  wire  _T_1899; 
  wire  _T_1900; 
  wire  _T_1911; 
  wire  _T_1913; 
  wire  _T_1914; 
  wire  _T_1919; 
  wire  _T_2049; 
  wire  _T_2059; 
  wire  _T_2061; 
  wire  _T_2062; 
  wire  _T_2067; 
  wire  _T_2081; 
  wire  _T_2099; 
  wire  _T_2101; 
  wire  _T_2102; 
  wire  _T_2103; 
  wire [5:0] _T_2108; 
  wire  _T_2109; 
  wire  _T_2110; 
  reg [5:0] _T_2112; 
  reg [31:0] _RAND_0;
  wire [5:0] _T_2114; 
  wire  _T_2115; 
  reg [2:0] _T_2123; 
  reg [31:0] _RAND_1;
  reg [2:0] _T_2124; 
  reg [31:0] _RAND_2;
  reg [3:0] _T_2125; 
  reg [31:0] _RAND_3;
  reg [5:0] _T_2126; 
  reg [31:0] _RAND_4;
  reg [31:0] _T_2127; 
  reg [31:0] _RAND_5;
  wire  _T_2128; 
  wire  _T_2129; 
  wire  _T_2130; 
  wire  _T_2132; 
  wire  _T_2133; 
  wire  _T_2134; 
  wire  _T_2136; 
  wire  _T_2137; 
  wire  _T_2138; 
  wire  _T_2140; 
  wire  _T_2141; 
  wire  _T_2142; 
  wire  _T_2144; 
  wire  _T_2145; 
  wire  _T_2146; 
  wire  _T_2148; 
  wire  _T_2149; 
  wire  _T_2151; 
  wire  _T_2152; 
  wire [22:0] _T_2154; 
  wire [7:0] _T_2155; 
  wire [7:0] _T_2156; 
  wire [5:0] _T_2157; 
  wire  _T_2158; 
  reg [5:0] _T_2160; 
  reg [31:0] _RAND_6;
  wire [5:0] _T_2162; 
  wire  _T_2163; 
  reg [2:0] _T_2171; 
  reg [31:0] _RAND_7;
  reg [1:0] _T_2172; 
  reg [31:0] _RAND_8;
  reg [3:0] _T_2173; 
  reg [31:0] _RAND_9;
  reg [5:0] _T_2174; 
  reg [31:0] _RAND_10;
  reg  _T_2175; 
  reg [31:0] _RAND_11;
  reg  _T_2176; 
  reg [31:0] _RAND_12;
  wire  _T_2177; 
  wire  _T_2178; 
  wire  _T_2179; 
  wire  _T_2181; 
  wire  _T_2182; 
  wire  _T_2183; 
  wire  _T_2185; 
  wire  _T_2186; 
  wire  _T_2187; 
  wire  _T_2189; 
  wire  _T_2190; 
  wire  _T_2191; 
  wire  _T_2193; 
  wire  _T_2194; 
  wire  _T_2195; 
  wire  _T_2197; 
  wire  _T_2198; 
  wire  _T_2199; 
  wire  _T_2201; 
  wire  _T_2202; 
  wire  _T_2204; 
  wire  _T_2254; 
  wire [5:0] _T_2259; 
  wire  _T_2260; 
  reg [5:0] _T_2262; 
  reg [31:0] _RAND_13;
  wire [5:0] _T_2264; 
  wire  _T_2265; 
  reg [2:0] _T_2273; 
  reg [31:0] _RAND_14;
  reg [2:0] _T_2274; 
  reg [31:0] _RAND_15;
  reg [3:0] _T_2275; 
  reg [31:0] _RAND_16;
  reg [5:0] _T_2276; 
  reg [31:0] _RAND_17;
  reg [31:0] _T_2277; 
  reg [31:0] _RAND_18;
  wire  _T_2278; 
  wire  _T_2279; 
  wire  _T_2280; 
  wire  _T_2282; 
  wire  _T_2283; 
  wire  _T_2284; 
  wire  _T_2286; 
  wire  _T_2287; 
  wire  _T_2288; 
  wire  _T_2290; 
  wire  _T_2291; 
  wire  _T_2292; 
  wire  _T_2294; 
  wire  _T_2295; 
  wire  _T_2296; 
  wire  _T_2298; 
  wire  _T_2299; 
  wire  _T_2301; 
  reg [63:0] _T_2302; 
  reg [63:0] _RAND_19;
  reg [5:0] _T_2312; 
  reg [31:0] _RAND_20;
  wire [5:0] _T_2314; 
  wire  _T_2315; 
  reg [5:0] _T_2331; 
  reg [31:0] _RAND_21;
  wire [5:0] _T_2333; 
  wire  _T_2334; 
  wire  _T_2344; 
  wire [63:0] _T_2346; 
  wire [63:0] _T_2347; 
  wire  _T_2348; 
  wire  _T_2349; 
  wire  _T_2351; 
  wire  _T_2352; 
  wire [63:0] _GEN_27; 
  wire  _T_2356; 
  wire  _T_2358; 
  wire  _T_2359; 
  wire [63:0] _T_2360; 
  wire [63:0] _T_2361; 
  wire [63:0] _T_2362; 
  wire  _T_2363; 
  wire  _T_2365; 
  wire  _T_2366; 
  wire [63:0] _GEN_28; 
  wire  _T_2367; 
  wire  _T_2368; 
  wire  _T_2369; 
  wire  _T_2370; 
  wire  _T_2372; 
  wire  _T_2373; 
  wire [63:0] _T_2374; 
  wire [63:0] _T_2375; 
  wire [63:0] _T_2376; 
  reg [31:0] _T_2377; 
  reg [31:0] _RAND_22;
  wire  _T_2378; 
  wire  _T_2379; 
  wire  _T_2380; 
  wire  _T_2381; 
  wire  _T_2382; 
  wire  _T_2383; 
  wire  _T_2385; 
  wire  _T_2386; 
  wire [31:0] _T_2388; 
  wire  _T_2391; 
  reg  _T_2392; 
  reg [31:0] _RAND_23;
  reg [5:0] _T_2401; 
  reg [31:0] _RAND_24;
  wire [5:0] _T_2403; 
  wire  _T_2404; 
  wire  _T_2414; 
  wire  _T_2415; 
  wire  _T_2416; 
  wire  _T_2417; 
  wire  _T_2418; 
  wire  _T_2419; 
  wire [1:0] _T_2420; 
  wire  _T_2421; 
  wire  _T_2423; 
  wire  _T_2425; 
  wire  _T_2426; 
  wire [1:0] _GEN_31; 
  wire  _T_2428; 
  wire [1:0] _T_2431; 
  wire  _T_2412; 
  wire  _T_2432; 
  wire  _T_2433; 
  wire  _T_2436; 
  wire  _T_2437; 
  wire [1:0] _GEN_32; 
  wire  _T_2438; 
  wire  _T_2427; 
  wire  _T_2439; 
  wire  _T_2440; 
  wire  _GEN_35; 
  wire  _GEN_49; 
  wire  _GEN_65; 
  wire  _GEN_75; 
  wire  _GEN_85; 
  wire  _GEN_95; 
  wire  _GEN_105; 
  wire  _GEN_115; 
  wire  _GEN_123; 
  wire  _GEN_133; 
  wire  _GEN_145; 
  wire  _GEN_157; 
  wire  _GEN_163; 
  wire  _GEN_169; 
  wire  _GEN_175; 
  wire  _GEN_187; 
  wire  _GEN_197; 
  wire  _GEN_211; 
  wire  _GEN_223; 
  wire  _GEN_233; 
  wire  _GEN_241; 
  dual_plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0)) plusarg_reader ( 
    .out(plusarg_reader_out)
  );
  assign _T_7 = io_in_a_bits_source[5:3]; 
  assign _T_8 = _T_7 == 3'h0; 
  assign _T_16 = _T_7 == 3'h1; 
  assign _T_24 = _T_7 == 3'h2; 
  assign _T_32 = _T_7 == 3'h3; 
  assign _T_40 = _T_7 == 3'h4; 
  assign _T_48 = _T_7 == 3'h5; 
  assign _T_56 = _T_7 == 3'h6; 
  assign _T_64 = _T_7 == 3'h7; 
  assign _T_70 = _T_8 | _T_16; 
  assign _T_71 = _T_70 | _T_24; 
  assign _T_72 = _T_71 | _T_32; 
  assign _T_73 = _T_72 | _T_40; 
  assign _T_74 = _T_73 | _T_48; 
  assign _T_75 = _T_74 | _T_56; 
  assign _T_76 = _T_75 | _T_64; 
  assign _T_78 = 23'hff << io_in_a_bits_size; 
  assign _T_79 = _T_78[7:0]; 
  assign _T_80 = ~ _T_79; 
  assign _GEN_33 = {{24'd0}, _T_80}; 
  assign _T_81 = io_in_a_bits_address & _GEN_33; 
  assign _T_82 = _T_81 == 32'h0; 
  assign _T_84 = io_in_a_bits_size[0]; 
  assign _T_85 = 2'h1 << _T_84; 
  assign _T_87 = _T_85 | 2'h1; 
  assign _T_88 = io_in_a_bits_size >= 4'h2; 
  assign _T_89 = _T_87[1]; 
  assign _T_90 = io_in_a_bits_address[1]; 
  assign _T_91 = _T_90 == 1'h0; 
  assign _T_93 = _T_89 & _T_91; 
  assign _T_94 = _T_88 | _T_93; 
  assign _T_96 = _T_89 & _T_90; 
  assign _T_97 = _T_88 | _T_96; 
  assign _T_98 = _T_87[0]; 
  assign _T_99 = io_in_a_bits_address[0]; 
  assign _T_100 = _T_99 == 1'h0; 
  assign _T_101 = _T_91 & _T_100; 
  assign _T_102 = _T_98 & _T_101; 
  assign _T_103 = _T_94 | _T_102; 
  assign _T_104 = _T_91 & _T_99; 
  assign _T_105 = _T_98 & _T_104; 
  assign _T_106 = _T_94 | _T_105; 
  assign _T_107 = _T_90 & _T_100; 
  assign _T_108 = _T_98 & _T_107; 
  assign _T_109 = _T_97 | _T_108; 
  assign _T_110 = _T_90 & _T_99; 
  assign _T_111 = _T_98 & _T_110; 
  assign _T_112 = _T_97 | _T_111; 
  assign _T_115 = {_T_112,_T_109,_T_106,_T_103}; 
  assign _T_246 = io_in_a_bits_opcode == 3'h6; 
  assign _T_248 = io_in_a_bits_address ^ 32'h80000000; 
  assign _T_249 = {1'b0,$signed(_T_248)}; 
  assign _T_250 = $signed(_T_249) & $signed(-33'sh80000000); 
  assign _T_251 = $signed(_T_250); 
  assign _T_252 = $signed(_T_251) == $signed(33'sh0); 
  assign _T_253 = io_in_a_bits_address ^ 32'h40000000; 
  assign _T_254 = {1'b0,$signed(_T_253)}; 
  assign _T_255 = $signed(_T_254) & $signed(-33'sh20000000); 
  assign _T_256 = $signed(_T_255); 
  assign _T_257 = $signed(_T_256) == $signed(33'sh0); 
  assign _T_258 = _T_252 | _T_257; 
  assign _T_261 = io_in_a_bits_size <= 4'h6; 
  assign _T_264 = io_in_a_bits_address ^ 32'h10000000; 
  assign _T_265 = {1'b0,$signed(_T_264)}; 
  assign _T_266 = $signed(_T_265) & $signed(-33'sh10000000); 
  assign _T_267 = $signed(_T_266); 
  assign _T_268 = $signed(_T_267) == $signed(33'sh0); 
  assign _T_269 = _T_261 & _T_268; 
  assign _T_273 = _T_269 | reset; 
  assign _T_274 = _T_273 == 1'h0; 
  assign _T_343 = _T_8 ? _T_261 : 1'h0; 
  assign _T_360 = _T_343 | reset; 
  assign _T_361 = _T_360 == 1'h0; 
  assign _T_363 = _T_76 | reset; 
  assign _T_364 = _T_363 == 1'h0; 
  assign _T_367 = _T_88 | reset; 
  assign _T_368 = _T_367 == 1'h0; 
  assign _T_370 = _T_82 | reset; 
  assign _T_371 = _T_370 == 1'h0; 
  assign _T_372 = io_in_a_bits_param <= 3'h2; 
  assign _T_374 = _T_372 | reset; 
  assign _T_375 = _T_374 == 1'h0; 
  assign _T_376 = ~ io_in_a_bits_mask; 
  assign _T_377 = _T_376 == 4'h0; 
  assign _T_379 = _T_377 | reset; 
  assign _T_380 = _T_379 == 1'h0; 
  assign _T_385 = io_in_a_bits_opcode == 3'h7; 
  assign _T_515 = io_in_a_bits_param != 3'h0; 
  assign _T_517 = _T_515 | reset; 
  assign _T_518 = _T_517 == 1'h0; 
  assign _T_528 = io_in_a_bits_opcode == 3'h4; 
  assign _T_549 = _T_258 | _T_268; 
  assign _T_550 = _T_261 & _T_549; 
  assign _T_553 = _T_550 | reset; 
  assign _T_554 = _T_553 == 1'h0; 
  assign _T_561 = io_in_a_bits_param == 3'h0; 
  assign _T_563 = _T_561 | reset; 
  assign _T_564 = _T_563 == 1'h0; 
  assign _T_565 = io_in_a_bits_mask == _T_115; 
  assign _T_567 = _T_565 | reset; 
  assign _T_568 = _T_567 == 1'h0; 
  assign _T_573 = io_in_a_bits_opcode == 3'h0; 
  assign _T_588 = _T_252 | _T_268; 
  assign _T_589 = _T_261 & _T_588; 
  assign _T_591 = io_in_a_bits_size <= 4'h8; 
  assign _T_599 = _T_591 & _T_257; 
  assign _T_601 = _T_589 | _T_599; 
  assign _T_603 = _T_601 | reset; 
  assign _T_604 = _T_603 == 1'h0; 
  assign _T_619 = io_in_a_bits_opcode == 3'h1; 
  assign _T_661 = ~ _T_115; 
  assign _T_662 = io_in_a_bits_mask & _T_661; 
  assign _T_663 = _T_662 == 4'h0; 
  assign _T_665 = _T_663 | reset; 
  assign _T_666 = _T_665 == 1'h0; 
  assign _T_667 = io_in_a_bits_opcode == 3'h2; 
  assign _T_669 = io_in_a_bits_size <= 4'h3; 
  assign _T_689 = _T_669 & _T_549; 
  assign _T_692 = _T_689 | reset; 
  assign _T_693 = _T_692 == 1'h0; 
  assign _T_700 = io_in_a_bits_param <= 3'h4; 
  assign _T_702 = _T_700 | reset; 
  assign _T_703 = _T_702 == 1'h0; 
  assign _T_708 = io_in_a_bits_opcode == 3'h3; 
  assign _T_741 = io_in_a_bits_param <= 3'h3; 
  assign _T_743 = _T_741 | reset; 
  assign _T_744 = _T_743 == 1'h0; 
  assign _T_749 = io_in_a_bits_opcode == 3'h5; 
  assign _T_795 = io_in_d_bits_opcode <= 3'h6; 
  assign _T_797 = _T_795 | reset; 
  assign _T_798 = _T_797 == 1'h0; 
  assign _T_801 = io_in_d_bits_source[5:3]; 
  assign _T_802 = _T_801 == 3'h0; 
  assign _T_810 = _T_801 == 3'h1; 
  assign _T_818 = _T_801 == 3'h2; 
  assign _T_826 = _T_801 == 3'h3; 
  assign _T_834 = _T_801 == 3'h4; 
  assign _T_842 = _T_801 == 3'h5; 
  assign _T_850 = _T_801 == 3'h6; 
  assign _T_858 = _T_801 == 3'h7; 
  assign _T_864 = _T_802 | _T_810; 
  assign _T_865 = _T_864 | _T_818; 
  assign _T_866 = _T_865 | _T_826; 
  assign _T_867 = _T_866 | _T_834; 
  assign _T_868 = _T_867 | _T_842; 
  assign _T_869 = _T_868 | _T_850; 
  assign _T_870 = _T_869 | _T_858; 
  assign _T_871 = io_in_d_bits_sink < 1'h1; 
  assign _T_872 = io_in_d_bits_opcode == 3'h6; 
  assign _T_874 = _T_870 | reset; 
  assign _T_875 = _T_874 == 1'h0; 
  assign _T_876 = io_in_d_bits_size >= 4'h2; 
  assign _T_878 = _T_876 | reset; 
  assign _T_879 = _T_878 == 1'h0; 
  assign _T_880 = io_in_d_bits_param == 2'h0; 
  assign _T_882 = _T_880 | reset; 
  assign _T_883 = _T_882 == 1'h0; 
  assign _T_884 = io_in_d_bits_corrupt == 1'h0; 
  assign _T_886 = _T_884 | reset; 
  assign _T_887 = _T_886 == 1'h0; 
  assign _T_888 = io_in_d_bits_denied == 1'h0; 
  assign _T_890 = _T_888 | reset; 
  assign _T_891 = _T_890 == 1'h0; 
  assign _T_892 = io_in_d_bits_opcode == 3'h4; 
  assign _T_897 = _T_871 | reset; 
  assign _T_898 = _T_897 == 1'h0; 
  assign _T_903 = io_in_d_bits_param <= 2'h2; 
  assign _T_905 = _T_903 | reset; 
  assign _T_906 = _T_905 == 1'h0; 
  assign _T_907 = io_in_d_bits_param != 2'h2; 
  assign _T_909 = _T_907 | reset; 
  assign _T_910 = _T_909 == 1'h0; 
  assign _T_920 = io_in_d_bits_opcode == 3'h5; 
  assign _T_940 = _T_888 | io_in_d_bits_corrupt; 
  assign _T_942 = _T_940 | reset; 
  assign _T_943 = _T_942 == 1'h0; 
  assign _T_949 = io_in_d_bits_opcode == 3'h0; 
  assign _T_966 = io_in_d_bits_opcode == 3'h1; 
  assign _T_984 = io_in_d_bits_opcode == 3'h2; 
  assign _T_1521 = io_in_c_bits_source[5:3]; 
  assign _T_1522 = _T_1521 == 3'h0; 
  assign _T_1530 = _T_1521 == 3'h1; 
  assign _T_1538 = _T_1521 == 3'h2; 
  assign _T_1546 = _T_1521 == 3'h3; 
  assign _T_1554 = _T_1521 == 3'h4; 
  assign _T_1562 = _T_1521 == 3'h5; 
  assign _T_1570 = _T_1521 == 3'h6; 
  assign _T_1578 = _T_1521 == 3'h7; 
  assign _T_1584 = _T_1522 | _T_1530; 
  assign _T_1585 = _T_1584 | _T_1538; 
  assign _T_1586 = _T_1585 | _T_1546; 
  assign _T_1587 = _T_1586 | _T_1554; 
  assign _T_1588 = _T_1587 | _T_1562; 
  assign _T_1589 = _T_1588 | _T_1570; 
  assign _T_1590 = _T_1589 | _T_1578; 
  assign _T_1592 = 23'hff << io_in_c_bits_size; 
  assign _T_1593 = _T_1592[7:0]; 
  assign _T_1594 = ~ _T_1593; 
  assign _GEN_34 = {{24'd0}, _T_1594}; 
  assign _T_1595 = io_in_c_bits_address & _GEN_34; 
  assign _T_1596 = _T_1595 == 32'h0; 
  assign _T_1597 = io_in_c_bits_address ^ 32'h80000000; 
  assign _T_1598 = {1'b0,$signed(_T_1597)}; 
  assign _T_1599 = $signed(_T_1598) & $signed(-33'sh80000000); 
  assign _T_1600 = $signed(_T_1599); 
  assign _T_1601 = $signed(_T_1600) == $signed(33'sh0); 
  assign _T_1602 = io_in_c_bits_address ^ 32'h40000000; 
  assign _T_1603 = {1'b0,$signed(_T_1602)}; 
  assign _T_1604 = $signed(_T_1603) & $signed(-33'sh20000000); 
  assign _T_1605 = $signed(_T_1604); 
  assign _T_1606 = $signed(_T_1605) == $signed(33'sh0); 
  assign _T_1607 = io_in_c_bits_address ^ 32'h10000000; 
  assign _T_1608 = {1'b0,$signed(_T_1607)}; 
  assign _T_1609 = $signed(_T_1608) & $signed(-33'sh10000000); 
  assign _T_1610 = $signed(_T_1609); 
  assign _T_1611 = $signed(_T_1610) == $signed(33'sh0); 
  assign _T_1613 = _T_1601 | _T_1606; 
  assign _T_1614 = _T_1613 | _T_1611; 
  assign _T_1745 = io_in_c_bits_opcode == 3'h4; 
  assign _T_1747 = _T_1614 | reset; 
  assign _T_1748 = _T_1747 == 1'h0; 
  assign _T_1750 = _T_1590 | reset; 
  assign _T_1751 = _T_1750 == 1'h0; 
  assign _T_1752 = io_in_c_bits_size >= 4'h2; 
  assign _T_1754 = _T_1752 | reset; 
  assign _T_1755 = _T_1754 == 1'h0; 
  assign _T_1757 = _T_1596 | reset; 
  assign _T_1758 = _T_1757 == 1'h0; 
  assign _T_1759 = io_in_c_bits_param <= 3'h5; 
  assign _T_1761 = _T_1759 | reset; 
  assign _T_1762 = _T_1761 == 1'h0; 
  assign _T_1763 = io_in_c_bits_corrupt == 1'h0; 
  assign _T_1765 = _T_1763 | reset; 
  assign _T_1766 = _T_1765 == 1'h0; 
  assign _T_1767 = io_in_c_bits_opcode == 3'h5; 
  assign _T_1785 = io_in_c_bits_opcode == 3'h6; 
  assign _T_1800 = io_in_c_bits_size <= 4'h6; 
  assign _T_1808 = _T_1800 & _T_1611; 
  assign _T_1812 = _T_1808 | reset; 
  assign _T_1813 = _T_1812 == 1'h0; 
  assign _T_1882 = _T_1522 ? _T_1800 : 1'h0; 
  assign _T_1899 = _T_1882 | reset; 
  assign _T_1900 = _T_1899 == 1'h0; 
  assign _T_1911 = io_in_c_bits_param <= 3'h2; 
  assign _T_1913 = _T_1911 | reset; 
  assign _T_1914 = _T_1913 == 1'h0; 
  assign _T_1919 = io_in_c_bits_opcode == 3'h7; 
  assign _T_2049 = io_in_c_bits_opcode == 3'h0; 
  assign _T_2059 = io_in_c_bits_param == 3'h0; 
  assign _T_2061 = _T_2059 | reset; 
  assign _T_2062 = _T_2061 == 1'h0; 
  assign _T_2067 = io_in_c_bits_opcode == 3'h1; 
  assign _T_2081 = io_in_c_bits_opcode == 3'h2; 
  assign _T_2099 = io_in_e_bits_sink < 1'h1; 
  assign _T_2101 = _T_2099 | reset; 
  assign _T_2102 = _T_2101 == 1'h0; 
  assign _T_2103 = io_in_a_ready & io_in_a_valid; 
  assign _T_2108 = _T_80[7:2]; 
  assign _T_2109 = io_in_a_bits_opcode[2]; 
  assign _T_2110 = _T_2109 == 1'h0; 
  assign _T_2114 = _T_2112 - 6'h1; 
  assign _T_2115 = _T_2112 == 6'h0; 
  assign _T_2128 = _T_2115 == 1'h0; 
  assign _T_2129 = io_in_a_valid & _T_2128; 
  assign _T_2130 = io_in_a_bits_opcode == _T_2123; 
  assign _T_2132 = _T_2130 | reset; 
  assign _T_2133 = _T_2132 == 1'h0; 
  assign _T_2134 = io_in_a_bits_param == _T_2124; 
  assign _T_2136 = _T_2134 | reset; 
  assign _T_2137 = _T_2136 == 1'h0; 
  assign _T_2138 = io_in_a_bits_size == _T_2125; 
  assign _T_2140 = _T_2138 | reset; 
  assign _T_2141 = _T_2140 == 1'h0; 
  assign _T_2142 = io_in_a_bits_source == _T_2126; 
  assign _T_2144 = _T_2142 | reset; 
  assign _T_2145 = _T_2144 == 1'h0; 
  assign _T_2146 = io_in_a_bits_address == _T_2127; 
  assign _T_2148 = _T_2146 | reset; 
  assign _T_2149 = _T_2148 == 1'h0; 
  assign _T_2151 = _T_2103 & _T_2115; 
  assign _T_2152 = io_in_d_ready & io_in_d_valid; 
  assign _T_2154 = 23'hff << io_in_d_bits_size; 
  assign _T_2155 = _T_2154[7:0]; 
  assign _T_2156 = ~ _T_2155; 
  assign _T_2157 = _T_2156[7:2]; 
  assign _T_2158 = io_in_d_bits_opcode[0]; 
  assign _T_2162 = _T_2160 - 6'h1; 
  assign _T_2163 = _T_2160 == 6'h0; 
  assign _T_2177 = _T_2163 == 1'h0; 
  assign _T_2178 = io_in_d_valid & _T_2177; 
  assign _T_2179 = io_in_d_bits_opcode == _T_2171; 
  assign _T_2181 = _T_2179 | reset; 
  assign _T_2182 = _T_2181 == 1'h0; 
  assign _T_2183 = io_in_d_bits_param == _T_2172; 
  assign _T_2185 = _T_2183 | reset; 
  assign _T_2186 = _T_2185 == 1'h0; 
  assign _T_2187 = io_in_d_bits_size == _T_2173; 
  assign _T_2189 = _T_2187 | reset; 
  assign _T_2190 = _T_2189 == 1'h0; 
  assign _T_2191 = io_in_d_bits_source == _T_2174; 
  assign _T_2193 = _T_2191 | reset; 
  assign _T_2194 = _T_2193 == 1'h0; 
  assign _T_2195 = io_in_d_bits_sink == _T_2175; 
  assign _T_2197 = _T_2195 | reset; 
  assign _T_2198 = _T_2197 == 1'h0; 
  assign _T_2199 = io_in_d_bits_denied == _T_2176; 
  assign _T_2201 = _T_2199 | reset; 
  assign _T_2202 = _T_2201 == 1'h0; 
  assign _T_2204 = _T_2152 & _T_2163; 
  assign _T_2254 = io_in_c_ready & io_in_c_valid; 
  assign _T_2259 = _T_1594[7:2]; 
  assign _T_2260 = io_in_c_bits_opcode[0]; 
  assign _T_2264 = _T_2262 - 6'h1; 
  assign _T_2265 = _T_2262 == 6'h0; 
  assign _T_2278 = _T_2265 == 1'h0; 
  assign _T_2279 = io_in_c_valid & _T_2278; 
  assign _T_2280 = io_in_c_bits_opcode == _T_2273; 
  assign _T_2282 = _T_2280 | reset; 
  assign _T_2283 = _T_2282 == 1'h0; 
  assign _T_2284 = io_in_c_bits_param == _T_2274; 
  assign _T_2286 = _T_2284 | reset; 
  assign _T_2287 = _T_2286 == 1'h0; 
  assign _T_2288 = io_in_c_bits_size == _T_2275; 
  assign _T_2290 = _T_2288 | reset; 
  assign _T_2291 = _T_2290 == 1'h0; 
  assign _T_2292 = io_in_c_bits_source == _T_2276; 
  assign _T_2294 = _T_2292 | reset; 
  assign _T_2295 = _T_2294 == 1'h0; 
  assign _T_2296 = io_in_c_bits_address == _T_2277; 
  assign _T_2298 = _T_2296 | reset; 
  assign _T_2299 = _T_2298 == 1'h0; 
  assign _T_2301 = _T_2254 & _T_2265; 
  assign _T_2314 = _T_2312 - 6'h1; 
  assign _T_2315 = _T_2312 == 6'h0; 
  assign _T_2333 = _T_2331 - 6'h1; 
  assign _T_2334 = _T_2331 == 6'h0; 
  assign _T_2344 = _T_2103 & _T_2315; 
  assign _T_2346 = 64'h1 << io_in_a_bits_source; 
  assign _T_2347 = _T_2302 >> io_in_a_bits_source; 
  assign _T_2348 = _T_2347[0]; 
  assign _T_2349 = _T_2348 == 1'h0; 
  assign _T_2351 = _T_2349 | reset; 
  assign _T_2352 = _T_2351 == 1'h0; 
  assign _GEN_27 = _T_2344 ? _T_2346 : 64'h0; 
  assign _T_2356 = _T_2152 & _T_2334; 
  assign _T_2358 = _T_872 == 1'h0; 
  assign _T_2359 = _T_2356 & _T_2358; 
  assign _T_2360 = 64'h1 << io_in_d_bits_source; 
  assign _T_2361 = _GEN_27 | _T_2302; 
  assign _T_2362 = _T_2361 >> io_in_d_bits_source; 
  assign _T_2363 = _T_2362[0]; 
  assign _T_2365 = _T_2363 | reset; 
  assign _T_2366 = _T_2365 == 1'h0; 
  assign _GEN_28 = _T_2359 ? _T_2360 : 64'h0; 
  assign _T_2367 = _GEN_27 != _GEN_28; 
  assign _T_2368 = _GEN_27 != 64'h0; 
  assign _T_2369 = _T_2368 == 1'h0; 
  assign _T_2370 = _T_2367 | _T_2369; 
  assign _T_2372 = _T_2370 | reset; 
  assign _T_2373 = _T_2372 == 1'h0; 
  assign _T_2374 = _T_2302 | _GEN_27; 
  assign _T_2375 = ~ _GEN_28; 
  assign _T_2376 = _T_2374 & _T_2375; 
  assign _T_2378 = _T_2302 != 64'h0; 
  assign _T_2379 = _T_2378 == 1'h0; 
  assign _T_2380 = plusarg_reader_out == 32'h0; 
  assign _T_2381 = _T_2379 | _T_2380; 
  assign _T_2382 = _T_2377 < plusarg_reader_out; 
  assign _T_2383 = _T_2381 | _T_2382; 
  assign _T_2385 = _T_2383 | reset; 
  assign _T_2386 = _T_2385 == 1'h0; 
  assign _T_2388 = _T_2377 + 32'h1; 
  assign _T_2391 = _T_2103 | _T_2152; 
  assign _T_2403 = _T_2401 - 6'h1; 
  assign _T_2404 = _T_2401 == 6'h0; 
  assign _T_2414 = _T_2152 & _T_2404; 
  assign _T_2415 = io_in_d_bits_opcode[2]; 
  assign _T_2416 = io_in_d_bits_opcode[1]; 
  assign _T_2417 = _T_2416 == 1'h0; 
  assign _T_2418 = _T_2415 & _T_2417; 
  assign _T_2419 = _T_2414 & _T_2418; 
  assign _T_2420 = 2'h1 << io_in_d_bits_sink; 
  assign _T_2421 = _T_2392 >> io_in_d_bits_sink; 
  assign _T_2423 = _T_2421 == 1'h0; 
  assign _T_2425 = _T_2423 | reset; 
  assign _T_2426 = _T_2425 == 1'h0; 
  assign _GEN_31 = _T_2419 ? _T_2420 : 2'h0; 
  assign _T_2428 = io_in_e_ready & io_in_e_valid; 
  assign _T_2431 = 2'h1 << io_in_e_bits_sink; 
  assign _T_2412 = _GEN_31[0]; 
  assign _T_2432 = _T_2412 | _T_2392; 
  assign _T_2433 = _T_2432 >> io_in_e_bits_sink; 
  assign _T_2436 = _T_2433 | reset; 
  assign _T_2437 = _T_2436 == 1'h0; 
  assign _GEN_32 = _T_2428 ? _T_2431 : 2'h0; 
  assign _T_2438 = _T_2392 | _T_2412; 
  assign _T_2427 = _GEN_32[0]; 
  assign _T_2439 = ~ _T_2427; 
  assign _T_2440 = _T_2438 & _T_2439; 
  assign _GEN_35 = io_in_a_valid & _T_246; 
  assign _GEN_49 = io_in_a_valid & _T_385; 
  assign _GEN_65 = io_in_a_valid & _T_528; 
  assign _GEN_75 = io_in_a_valid & _T_573; 
  assign _GEN_85 = io_in_a_valid & _T_619; 
  assign _GEN_95 = io_in_a_valid & _T_667; 
  assign _GEN_105 = io_in_a_valid & _T_708; 
  assign _GEN_115 = io_in_a_valid & _T_749; 
  assign _GEN_123 = io_in_d_valid & _T_872; 
  assign _GEN_133 = io_in_d_valid & _T_892; 
  assign _GEN_145 = io_in_d_valid & _T_920; 
  assign _GEN_157 = io_in_d_valid & _T_949; 
  assign _GEN_163 = io_in_d_valid & _T_966; 
  assign _GEN_169 = io_in_d_valid & _T_984; 
  assign _GEN_175 = io_in_c_valid & _T_1745; 
  assign _GEN_187 = io_in_c_valid & _T_1767; 
  assign _GEN_197 = io_in_c_valid & _T_1785; 
  assign _GEN_211 = io_in_c_valid & _T_1919; 
  assign _GEN_223 = io_in_c_valid & _T_2049; 
  assign _GEN_233 = io_in_c_valid & _T_2067; 
  assign _GEN_241 = io_in_c_valid & _T_2081; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2112 = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_2123 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2124 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_2125 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_2126 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_2127 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_2160 = _RAND_6[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_2171 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_2172 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_2173 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_2174 = _RAND_10[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_2175 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_2176 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_2262 = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_2273 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_2274 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_2275 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_2276 = _RAND_17[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_2277 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  _T_2302 = _RAND_19[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_2312 = _RAND_20[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_2331 = _RAND_21[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_2377 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_2392 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_2401 = _RAND_24[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_2112 <= 6'h0;
    end else begin
      if (_T_2103) begin
        if (_T_2115) begin
          if (_T_2110) begin
            _T_2112 <= _T_2108;
          end else begin
            _T_2112 <= 6'h0;
          end
        end else begin
          _T_2112 <= _T_2114;
        end
      end
    end
    if (_T_2151) begin
      _T_2123 <= io_in_a_bits_opcode;
    end
    if (_T_2151) begin
      _T_2124 <= io_in_a_bits_param;
    end
    if (_T_2151) begin
      _T_2125 <= io_in_a_bits_size;
    end
    if (_T_2151) begin
      _T_2126 <= io_in_a_bits_source;
    end
    if (_T_2151) begin
      _T_2127 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_2160 <= 6'h0;
    end else begin
      if (_T_2152) begin
        if (_T_2163) begin
          if (_T_2158) begin
            _T_2160 <= _T_2157;
          end else begin
            _T_2160 <= 6'h0;
          end
        end else begin
          _T_2160 <= _T_2162;
        end
      end
    end
    if (_T_2204) begin
      _T_2171 <= io_in_d_bits_opcode;
    end
    if (_T_2204) begin
      _T_2172 <= io_in_d_bits_param;
    end
    if (_T_2204) begin
      _T_2173 <= io_in_d_bits_size;
    end
    if (_T_2204) begin
      _T_2174 <= io_in_d_bits_source;
    end
    if (_T_2204) begin
      _T_2175 <= io_in_d_bits_sink;
    end
    if (_T_2204) begin
      _T_2176 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_2262 <= 6'h0;
    end else begin
      if (_T_2254) begin
        if (_T_2265) begin
          if (_T_2260) begin
            _T_2262 <= _T_2259;
          end else begin
            _T_2262 <= 6'h0;
          end
        end else begin
          _T_2262 <= _T_2264;
        end
      end
    end
    if (_T_2301) begin
      _T_2273 <= io_in_c_bits_opcode;
    end
    if (_T_2301) begin
      _T_2274 <= io_in_c_bits_param;
    end
    if (_T_2301) begin
      _T_2275 <= io_in_c_bits_size;
    end
    if (_T_2301) begin
      _T_2276 <= io_in_c_bits_source;
    end
    if (_T_2301) begin
      _T_2277 <= io_in_c_bits_address;
    end
    if (reset) begin
      _T_2302 <= 64'h0;
    end else begin
      _T_2302 <= _T_2376;
    end
    if (reset) begin
      _T_2312 <= 6'h0;
    end else begin
      if (_T_2103) begin
        if (_T_2315) begin
          if (_T_2110) begin
            _T_2312 <= _T_2108;
          end else begin
            _T_2312 <= 6'h0;
          end
        end else begin
          _T_2312 <= _T_2314;
        end
      end
    end
    if (reset) begin
      _T_2331 <= 6'h0;
    end else begin
      if (_T_2152) begin
        if (_T_2334) begin
          if (_T_2158) begin
            _T_2331 <= _T_2157;
          end else begin
            _T_2331 <= 6'h0;
          end
        end else begin
          _T_2331 <= _T_2333;
        end
      end
    end
    if (reset) begin
      _T_2377 <= 32'h0;
    end else begin
      if (_T_2391) begin
        _T_2377 <= 32'h0;
      end else begin
        _T_2377 <= _T_2388;
      end
    end
    if (reset) begin
      _T_2392 <= 1'h0;
    end else begin
      _T_2392 <= _T_2440;
    end
    if (reset) begin
      _T_2401 <= 6'h0;
    end else begin
      if (_T_2152) begin
        if (_T_2404) begin
          if (_T_2158) begin
            _T_2401 <= _T_2157;
          end else begin
            _T_2401 <= 6'h0;
          end
        end else begin
          _T_2401 <= _T_2403;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel has invalid opcode (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:39 assert (TLMessages.isA(bundle.opcode), \"'A' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:46 assert (visible(edge.address(bundle), bundle.source, edge), \"'A' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_274) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_274) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_361) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_361) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_364) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_364) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_368) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_368) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_371) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_371) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_375) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_375) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_380) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_380) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:56 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_274) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_274) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_361) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_361) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_364) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_364) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_368) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_368) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_371) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_371) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_375) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_375) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_518) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_518) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_380) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_380) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:68 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_554) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_554) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_364) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_364) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_371) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_371) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_564) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_564) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_568) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_568) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:77 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_604) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_604) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_364) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_364) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_371) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_371) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_564) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_564) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_568) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_568) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_604) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_604) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_364) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_364) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_371) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_371) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_564) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_564) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_666) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_666) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_693) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_693) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_364) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_364) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_371) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_371) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_703) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_703) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_568) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_568) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_693) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_693) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_364) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_364) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_371) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_371) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_744) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_744) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_568) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_568) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_604) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_604) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_364) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_364) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_371) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_371) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_568) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_568) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:117 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_798) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_798) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_875) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_875) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_879) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_879) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_883) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_883) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_887) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_887) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_891) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_891) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_875) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_875) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_898) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:285 assert (sink_ok, \"'D' channel Grant carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_898) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_879) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_879) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_906) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_906) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_910) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_910) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_887) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_887) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is denied (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:290 assert (deny_put_ok || !bundle.denied, \"'D' channel Grant is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_875) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_875) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_898) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:295 assert (sink_ok, \"'D' channel GrantData carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_898) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_879) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_879) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_906) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_906) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_910) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_910) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_943) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_943) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:300 assert (deny_get_ok || !bundle.denied, \"'D' channel GrantData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_157 & _T_875) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_157 & _T_875) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_157 & _T_883) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_157 & _T_883) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_157 & _T_887) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_157 & _T_887) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is denied (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:308 assert (deny_put_ok || !bundle.denied, \"'D' channel AccessAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_875) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_875) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_883) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_883) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_943) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_943) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:316 assert (deny_get_ok || !bundle.denied, \"'D' channel AccessAckData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_169 & _T_875) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_169 & _T_875) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_169 & _T_883) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_169 & _T_883) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_169 & _T_887) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_169 & _T_887) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is denied (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:324 assert (deny_put_ok || !bundle.denied, \"'D' channel HintAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel has invalid opcode (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:122 assert (TLMessages.isB(bundle.opcode), \"'B' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:124 assert (visible(edge.address(bundle), bundle.source, edge), \"'B' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Probe type unsupported by client (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:133 assert (edge.client.supportsProbe(bundle.source, bundle.size), \"'B' channel carries Probe type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:134 assert (address_ok, \"'B' channel Probe carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries source that is not first source (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:135 assert (legal_source, \"'B' channel Probe carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:136 assert (is_aligned, \"'B' channel Probe address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:137 assert (TLPermissions.isCap(bundle.param), \"'B' channel Probe carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe contains invalid mask (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:138 assert (bundle.mask === mask, \"'B' channel Probe contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe is corrupt (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:139 assert (!bundle.corrupt, \"'B' channel Probe is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Get type unsupported by client (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:143 assert (edge.client.supportsGet(bundle.source, bundle.size), \"'B' channel carries Get type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries unmanaged address (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:144 assert (address_ok, \"'B' channel Get carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries source that is not first source (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:145 assert (legal_source, \"'B' channel Get carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:146 assert (is_aligned, \"'B' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries invalid param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:147 assert (bundle.param === UInt(0), \"'B' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get contains invalid mask (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:148 assert (bundle.mask === mask, \"'B' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get is corrupt (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:149 assert (!bundle.corrupt, \"'B' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutFull type unsupported by client (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:153 assert (edge.client.supportsPutFull(bundle.source, bundle.size), \"'B' channel carries PutFull type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries unmanaged address (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:154 assert (address_ok, \"'B' channel PutFull carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries source that is not first source (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:155 assert (legal_source, \"'B' channel PutFull carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:156 assert (is_aligned, \"'B' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries invalid param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:157 assert (bundle.param === UInt(0), \"'B' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull contains invalid mask (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:158 assert (bundle.mask === mask, \"'B' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutPartial type unsupported by client (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:162 assert (edge.client.supportsPutPartial(bundle.source, bundle.size), \"'B' channel carries PutPartial type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:163 assert (address_ok, \"'B' channel PutPartial carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:164 assert (legal_source, \"'B' channel PutPartial carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:165 assert (is_aligned, \"'B' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries invalid param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:166 assert (bundle.param === UInt(0), \"'B' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial contains invalid mask (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:167 assert ((bundle.mask & ~mask) === UInt(0), \"'B' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Arithmetic type unsupported by client (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:171 assert (edge.client.supportsArithmetic(bundle.source, bundle.size), \"'B' channel carries Arithmetic type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:172 assert (address_ok, \"'B' channel Arithmetic carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:173 assert (legal_source, \"'B' channel Arithmetic carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:174 assert (is_aligned, \"'B' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries invalid opcode param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:175 assert (TLAtomics.isArithmetic(bundle.param), \"'B' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:176 assert (bundle.mask === mask, \"'B' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Logical type unsupported by client (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:180 assert (edge.client.supportsLogical(bundle.source, bundle.size), \"'B' channel carries Logical type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries unmanaged address (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:181 assert (address_ok, \"'B' channel Logical carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries source that is not first source (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:182 assert (legal_source, \"'B' channel Logical carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:183 assert (is_aligned, \"'B' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries invalid opcode param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:184 assert (TLAtomics.isLogical(bundle.param), \"'B' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical contains invalid mask (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:185 assert (bundle.mask === mask, \"'B' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Hint type unsupported by client (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:189 assert (edge.client.supportsHint(bundle.source, bundle.size), \"'B' channel carries Hint type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries unmanaged address (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:190 assert (address_ok, \"'B' channel Hint carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries source that is not first source (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:191 assert (legal_source, \"'B' channel Hint carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:192 assert (is_aligned, \"'B' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint contains invalid mask (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:193 assert (bundle.mask === mask, \"'B' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint is corrupt (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:194 assert (!bundle.corrupt, \"'B' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel has invalid opcode (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:199 assert (TLMessages.isC(bundle.opcode), \"'C' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:205 assert (visible(edge.address(bundle), bundle.source, edge), \"'C' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1748) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:208 assert (address_ok, \"'C' channel ProbeAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1748) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1751) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:209 assert (source_ok, \"'C' channel ProbeAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1751) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1755) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:210 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1755) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1758) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:211 assert (is_aligned, \"'C' channel ProbeAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1758) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1762) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:212 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAck carries invalid report param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1762) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1766) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck is corrupt (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:213 assert (!bundle.corrupt, \"'C' channel ProbeAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1766) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_187 & _T_1748) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:217 assert (address_ok, \"'C' channel ProbeAckData carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_187 & _T_1748) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_187 & _T_1751) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:218 assert (source_ok, \"'C' channel ProbeAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_187 & _T_1751) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_187 & _T_1755) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:219 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAckData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_187 & _T_1755) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_187 & _T_1758) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:220 assert (is_aligned, \"'C' channel ProbeAckData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_187 & _T_1758) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_187 & _T_1762) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:221 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAckData carries invalid report param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_187 & _T_1762) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1813) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:225 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries Release type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1813) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1900) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:226 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1900) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1751) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:227 assert (source_ok, \"'C' channel Release carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1751) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1755) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:228 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel Release smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1755) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1758) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:229 assert (is_aligned, \"'C' channel Release address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1758) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1914) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid shrink param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:230 assert (TLPermissions.isShrink(bundle.param), \"'C' channel Release carries invalid shrink param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1914) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_197 & _T_1766) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release is corrupt (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:231 assert (!bundle.corrupt, \"'C' channel Release is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_197 & _T_1766) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1813) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:235 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries ReleaseData type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1813) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1900) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:236 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1900) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1751) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:237 assert (source_ok, \"'C' channel ReleaseData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1751) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1755) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:238 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ReleaseData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1755) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1758) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:239 assert (is_aligned, \"'C' channel ReleaseData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1758) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_211 & _T_1914) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid shrink param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:240 assert (TLPermissions.isShrink(bundle.param), \"'C' channel ReleaseData carries invalid shrink param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_211 & _T_1914) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_1748) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:244 assert (address_ok, \"'C' channel AccessAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_1748) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_1751) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:245 assert (source_ok, \"'C' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_1751) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_1758) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:246 assert (is_aligned, \"'C' channel AccessAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_1758) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_2062) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:247 assert (bundle.param === UInt(0), \"'C' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_2062) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_1766) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck is corrupt (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:248 assert (!bundle.corrupt, \"'C' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_1766) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_1748) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:252 assert (address_ok, \"'C' channel AccessAckData carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_1748) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_1751) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:253 assert (source_ok, \"'C' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_1751) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_1758) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:254 assert (is_aligned, \"'C' channel AccessAckData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_1758) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_2062) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:255 assert (bundle.param === UInt(0), \"'C' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_2062) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1748) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:259 assert (address_ok, \"'C' channel HintAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1748) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1751) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:260 assert (source_ok, \"'C' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1751) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1758) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:261 assert (is_aligned, \"'C' channel HintAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1758) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_2062) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:262 assert (bundle.param === UInt(0), \"'C' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_2062) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1766) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck is corrupt (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:263 assert (!bundle.corrupt, \"'C' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1766) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_e_valid & _T_2102) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channels carries invalid sink ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:330 assert (sink_ok, \"'E' channels carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_e_valid & _T_2102) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2129 & _T_2133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2129 & _T_2133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2129 & _T_2137) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2129 & _T_2137) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2129 & _T_2141) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2129 & _T_2141) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2129 & _T_2145) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2129 & _T_2145) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2129 & _T_2149) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2129 & _T_2149) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2178 & _T_2182) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2178 & _T_2182) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2178 & _T_2186) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2178 & _T_2186) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2178 & _T_2190) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2178 & _T_2190) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2178 & _T_2194) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2178 & _T_2194) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2178 & _T_2198) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2178 & _T_2198) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2178 & _T_2202) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2178 & _T_2202) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:378 assert (b.bits.opcode === opcode, \"'B' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:379 assert (b.bits.param  === param,  \"'B' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel size changed within multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:380 assert (b.bits.size   === size,   \"'B' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel source changed within multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:381 assert (b.bits.source === source, \"'B' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:382 assert (b.bits.address=== address,\"'B' channel addresss changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2279 & _T_2283) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:401 assert (c.bits.opcode === opcode, \"'C' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2279 & _T_2283) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2279 & _T_2287) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:402 assert (c.bits.param  === param,  \"'C' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2279 & _T_2287) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2279 & _T_2291) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:403 assert (c.bits.size   === size,   \"'C' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2279 & _T_2291) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2279 & _T_2295) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:404 assert (c.bits.source === source, \"'C' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2279 & _T_2295) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2279 & _T_2299) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:405 assert (c.bits.address=== address,\"'C' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2279 & _T_2299) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2344 & _T_2352) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2344 & _T_2352) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2359 & _T_2366) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2359 & _T_2366) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2373) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2373) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2386) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:479 assert (!inflight.orR || limit === UInt(0) || watchdog < limit, \"TileLink timeout expired\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2386) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2419 & _T_2426) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:494 assert(!inflight(bundle.d.bits.sink), \"'D' channel re-used a sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2419 & _T_2426) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2428 & _T_2437) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at ChiplinkTest.scala:362:118)\n    at Monitor.scala:500 assert((d_set | inflight)(bundle.e.bits.sink), \"'E' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2428 & _T_2437) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLMonitor_18( 
  input         clock, 
  input         reset, 
  input         io_in_a_ready, 
  input         io_in_a_valid, 
  input  [2:0]  io_in_a_bits_opcode, 
  input  [2:0]  io_in_a_bits_param, 
  input  [2:0]  io_in_a_bits_size, 
  input  [6:0]  io_in_a_bits_source, 
  input  [28:0] io_in_a_bits_address, 
  input  [7:0]  io_in_a_bits_mask, 
  input         io_in_a_bits_corrupt, 
  input         io_in_c_ready, 
  input         io_in_c_valid, 
  input  [2:0]  io_in_c_bits_opcode, 
  input  [2:0]  io_in_c_bits_param, 
  input  [2:0]  io_in_c_bits_size, 
  input  [6:0]  io_in_c_bits_source, 
  input  [28:0] io_in_c_bits_address, 
  input         io_in_c_bits_corrupt, 
  input         io_in_d_ready, 
  input         io_in_d_valid, 
  input  [2:0]  io_in_d_bits_opcode, 
  input  [1:0]  io_in_d_bits_param, 
  input  [2:0]  io_in_d_bits_size, 
  input  [6:0]  io_in_d_bits_source, 
  input         io_in_d_bits_sink, 
  input         io_in_d_bits_denied, 
  input         io_in_d_bits_corrupt, 
  input         io_in_e_valid 
);
  wire [31:0] plusarg_reader_out; 
  wire [2:0] _T_7; 
  wire  _T_8; 
  wire  _T_16; 
  wire  _T_24; 
  wire  _T_32; 
  wire  _T_40; 
  wire  _T_48; 
  wire  _T_56; 
  wire  _T_64; 
  wire  _T_70; 
  wire  _T_71; 
  wire  _T_72; 
  wire  _T_73; 
  wire  _T_74; 
  wire  _T_75; 
  wire  _T_76; 
  wire [12:0] _T_78; 
  wire [5:0] _T_79; 
  wire [5:0] _T_80; 
  wire [28:0] _GEN_33; 
  wire [28:0] _T_81; 
  wire  _T_82; 
  wire [1:0] _T_84; 
  wire [3:0] _T_85; 
  wire [2:0] _T_86; 
  wire [2:0] _T_87; 
  wire  _T_88; 
  wire  _T_89; 
  wire  _T_90; 
  wire  _T_91; 
  wire  _T_93; 
  wire  _T_94; 
  wire  _T_96; 
  wire  _T_97; 
  wire  _T_98; 
  wire  _T_99; 
  wire  _T_100; 
  wire  _T_101; 
  wire  _T_102; 
  wire  _T_103; 
  wire  _T_104; 
  wire  _T_105; 
  wire  _T_106; 
  wire  _T_107; 
  wire  _T_108; 
  wire  _T_109; 
  wire  _T_110; 
  wire  _T_111; 
  wire  _T_112; 
  wire  _T_113; 
  wire  _T_114; 
  wire  _T_115; 
  wire  _T_116; 
  wire  _T_117; 
  wire  _T_118; 
  wire  _T_119; 
  wire  _T_120; 
  wire  _T_121; 
  wire  _T_122; 
  wire  _T_123; 
  wire  _T_124; 
  wire  _T_125; 
  wire  _T_126; 
  wire  _T_127; 
  wire  _T_128; 
  wire  _T_129; 
  wire  _T_130; 
  wire  _T_131; 
  wire  _T_132; 
  wire  _T_133; 
  wire  _T_134; 
  wire  _T_135; 
  wire  _T_136; 
  wire  _T_137; 
  wire  _T_138; 
  wire  _T_139; 
  wire [7:0] _T_146; 
  wire  _T_277; 
  wire  _T_279; 
  wire [28:0] _T_282; 
  wire [29:0] _T_283; 
  wire [29:0] _T_284; 
  wire [29:0] _T_285; 
  wire  _T_286; 
  wire  _T_287; 
  wire  _T_290; 
  wire  _T_291; 
  wire  _T_360; 
  wire  _T_377; 
  wire  _T_378; 
  wire  _T_380; 
  wire  _T_381; 
  wire  _T_384; 
  wire  _T_385; 
  wire  _T_387; 
  wire  _T_388; 
  wire  _T_389; 
  wire  _T_391; 
  wire  _T_392; 
  wire [7:0] _T_393; 
  wire  _T_394; 
  wire  _T_396; 
  wire  _T_397; 
  wire  _T_398; 
  wire  _T_400; 
  wire  _T_401; 
  wire  _T_402; 
  wire  _T_518; 
  wire  _T_520; 
  wire  _T_521; 
  wire  _T_531; 
  wire  _T_552; 
  wire  _T_554; 
  wire  _T_555; 
  wire  _T_556; 
  wire  _T_558; 
  wire  _T_559; 
  wire  _T_564; 
  wire  _T_593; 
  wire [7:0] _T_618; 
  wire [7:0] _T_619; 
  wire  _T_620; 
  wire  _T_622; 
  wire  _T_623; 
  wire  _T_624; 
  wire  _T_645; 
  wire  _T_647; 
  wire  _T_648; 
  wire  _T_653; 
  wire  _T_674; 
  wire  _T_676; 
  wire  _T_677; 
  wire  _T_682; 
  wire  _T_711; 
  wire  _T_713; 
  wire  _T_714; 
  wire [2:0] _T_717; 
  wire  _T_718; 
  wire  _T_726; 
  wire  _T_734; 
  wire  _T_742; 
  wire  _T_750; 
  wire  _T_758; 
  wire  _T_766; 
  wire  _T_774; 
  wire  _T_780; 
  wire  _T_781; 
  wire  _T_782; 
  wire  _T_783; 
  wire  _T_784; 
  wire  _T_785; 
  wire  _T_786; 
  wire  _T_787; 
  wire  _T_788; 
  wire  _T_790; 
  wire  _T_791; 
  wire  _T_792; 
  wire  _T_794; 
  wire  _T_795; 
  wire  _T_796; 
  wire  _T_798; 
  wire  _T_799; 
  wire  _T_800; 
  wire  _T_802; 
  wire  _T_803; 
  wire  _T_804; 
  wire  _T_806; 
  wire  _T_807; 
  wire  _T_808; 
  wire  _T_813; 
  wire  _T_814; 
  wire  _T_819; 
  wire  _T_821; 
  wire  _T_822; 
  wire  _T_823; 
  wire  _T_825; 
  wire  _T_826; 
  wire  _T_836; 
  wire  _T_856; 
  wire  _T_858; 
  wire  _T_859; 
  wire  _T_865; 
  wire  _T_882; 
  wire  _T_900; 
  wire [2:0] _T_1456; 
  wire  _T_1457; 
  wire  _T_1465; 
  wire  _T_1473; 
  wire  _T_1481; 
  wire  _T_1489; 
  wire  _T_1497; 
  wire  _T_1505; 
  wire  _T_1513; 
  wire  _T_1519; 
  wire  _T_1520; 
  wire  _T_1521; 
  wire  _T_1522; 
  wire  _T_1523; 
  wire  _T_1524; 
  wire  _T_1525; 
  wire [12:0] _T_1527; 
  wire [5:0] _T_1528; 
  wire [5:0] _T_1529; 
  wire [28:0] _GEN_34; 
  wire [28:0] _T_1530; 
  wire  _T_1531; 
  wire [28:0] _T_1532; 
  wire [29:0] _T_1533; 
  wire [29:0] _T_1534; 
  wire [29:0] _T_1535; 
  wire  _T_1536; 
  wire  _T_1668; 
  wire  _T_1670; 
  wire  _T_1671; 
  wire  _T_1673; 
  wire  _T_1674; 
  wire  _T_1675; 
  wire  _T_1677; 
  wire  _T_1678; 
  wire  _T_1680; 
  wire  _T_1681; 
  wire  _T_1682; 
  wire  _T_1684; 
  wire  _T_1685; 
  wire  _T_1686; 
  wire  _T_1688; 
  wire  _T_1689; 
  wire  _T_1690; 
  wire  _T_1708; 
  wire  _T_1710; 
  wire  _T_1718; 
  wire  _T_1721; 
  wire  _T_1722; 
  wire  _T_1791; 
  wire  _T_1808; 
  wire  _T_1809; 
  wire  _T_1820; 
  wire  _T_1822; 
  wire  _T_1823; 
  wire  _T_1828; 
  wire  _T_1944; 
  wire  _T_1954; 
  wire  _T_1956; 
  wire  _T_1957; 
  wire  _T_1962; 
  wire  _T_1976; 
  wire  _T_1998; 
  wire [2:0] _T_2003; 
  wire  _T_2004; 
  wire  _T_2005; 
  reg [2:0] _T_2007; 
  reg [31:0] _RAND_0;
  wire [2:0] _T_2009; 
  wire  _T_2010; 
  reg [2:0] _T_2018; 
  reg [31:0] _RAND_1;
  reg [2:0] _T_2019; 
  reg [31:0] _RAND_2;
  reg [2:0] _T_2020; 
  reg [31:0] _RAND_3;
  reg [6:0] _T_2021; 
  reg [31:0] _RAND_4;
  reg [28:0] _T_2022; 
  reg [31:0] _RAND_5;
  wire  _T_2023; 
  wire  _T_2024; 
  wire  _T_2025; 
  wire  _T_2027; 
  wire  _T_2028; 
  wire  _T_2029; 
  wire  _T_2031; 
  wire  _T_2032; 
  wire  _T_2033; 
  wire  _T_2035; 
  wire  _T_2036; 
  wire  _T_2037; 
  wire  _T_2039; 
  wire  _T_2040; 
  wire  _T_2041; 
  wire  _T_2043; 
  wire  _T_2044; 
  wire  _T_2046; 
  wire  _T_2047; 
  wire [12:0] _T_2049; 
  wire [5:0] _T_2050; 
  wire [5:0] _T_2051; 
  wire [2:0] _T_2052; 
  wire  _T_2053; 
  reg [2:0] _T_2055; 
  reg [31:0] _RAND_6;
  wire [2:0] _T_2057; 
  wire  _T_2058; 
  reg [2:0] _T_2066; 
  reg [31:0] _RAND_7;
  reg [1:0] _T_2067; 
  reg [31:0] _RAND_8;
  reg [2:0] _T_2068; 
  reg [31:0] _RAND_9;
  reg [6:0] _T_2069; 
  reg [31:0] _RAND_10;
  reg  _T_2070; 
  reg [31:0] _RAND_11;
  reg  _T_2071; 
  reg [31:0] _RAND_12;
  wire  _T_2072; 
  wire  _T_2073; 
  wire  _T_2074; 
  wire  _T_2076; 
  wire  _T_2077; 
  wire  _T_2078; 
  wire  _T_2080; 
  wire  _T_2081; 
  wire  _T_2082; 
  wire  _T_2084; 
  wire  _T_2085; 
  wire  _T_2086; 
  wire  _T_2088; 
  wire  _T_2089; 
  wire  _T_2090; 
  wire  _T_2092; 
  wire  _T_2093; 
  wire  _T_2094; 
  wire  _T_2096; 
  wire  _T_2097; 
  wire  _T_2099; 
  wire  _T_2149; 
  wire [2:0] _T_2154; 
  wire  _T_2155; 
  reg [2:0] _T_2157; 
  reg [31:0] _RAND_13;
  wire [2:0] _T_2159; 
  wire  _T_2160; 
  reg [2:0] _T_2168; 
  reg [31:0] _RAND_14;
  reg [2:0] _T_2169; 
  reg [31:0] _RAND_15;
  reg [2:0] _T_2170; 
  reg [31:0] _RAND_16;
  reg [6:0] _T_2171; 
  reg [31:0] _RAND_17;
  reg [28:0] _T_2172; 
  reg [31:0] _RAND_18;
  wire  _T_2173; 
  wire  _T_2174; 
  wire  _T_2175; 
  wire  _T_2177; 
  wire  _T_2178; 
  wire  _T_2179; 
  wire  _T_2181; 
  wire  _T_2182; 
  wire  _T_2183; 
  wire  _T_2185; 
  wire  _T_2186; 
  wire  _T_2187; 
  wire  _T_2189; 
  wire  _T_2190; 
  wire  _T_2191; 
  wire  _T_2193; 
  wire  _T_2194; 
  wire  _T_2196; 
  reg [127:0] _T_2197; 
  reg [127:0] _RAND_19;
  reg [2:0] _T_2207; 
  reg [31:0] _RAND_20;
  wire [2:0] _T_2209; 
  wire  _T_2210; 
  reg [2:0] _T_2226; 
  reg [31:0] _RAND_21;
  wire [2:0] _T_2228; 
  wire  _T_2229; 
  wire  _T_2239; 
  wire [127:0] _T_2241; 
  wire [127:0] _T_2242; 
  wire  _T_2243; 
  wire  _T_2244; 
  wire  _T_2246; 
  wire  _T_2247; 
  wire [127:0] _GEN_27; 
  wire  _T_2251; 
  wire  _T_2253; 
  wire  _T_2254; 
  wire [127:0] _T_2255; 
  wire [127:0] _T_2256; 
  wire [127:0] _T_2257; 
  wire  _T_2258; 
  wire  _T_2260; 
  wire  _T_2261; 
  wire [127:0] _GEN_28; 
  wire  _T_2262; 
  wire  _T_2263; 
  wire  _T_2264; 
  wire  _T_2265; 
  wire  _T_2267; 
  wire  _T_2268; 
  wire [127:0] _T_2269; 
  wire [127:0] _T_2270; 
  wire [127:0] _T_2271; 
  reg [31:0] _T_2272; 
  reg [31:0] _RAND_22;
  wire  _T_2273; 
  wire  _T_2274; 
  wire  _T_2275; 
  wire  _T_2276; 
  wire  _T_2277; 
  wire  _T_2278; 
  wire  _T_2280; 
  wire  _T_2281; 
  wire [31:0] _T_2283; 
  wire  _T_2286; 
  reg  _T_2287; 
  reg [31:0] _RAND_23;
  reg [2:0] _T_2296; 
  reg [31:0] _RAND_24;
  wire [2:0] _T_2298; 
  wire  _T_2299; 
  wire  _T_2309; 
  wire  _T_2310; 
  wire  _T_2311; 
  wire  _T_2312; 
  wire  _T_2313; 
  wire  _T_2314; 
  wire [1:0] _T_2315; 
  wire  _T_2316; 
  wire  _T_2318; 
  wire  _T_2320; 
  wire  _T_2321; 
  wire [1:0] _GEN_31; 
  wire  _T_2307; 
  wire  _T_2327; 
  wire  _T_2331; 
  wire  _T_2332; 
  wire [1:0] _GEN_32; 
  wire  _T_2333; 
  wire  _T_2322; 
  wire  _T_2334; 
  wire  _T_2335; 
  wire  _GEN_35; 
  wire  _GEN_51; 
  wire  _GEN_69; 
  wire  _GEN_81; 
  wire  _GEN_91; 
  wire  _GEN_101; 
  wire  _GEN_111; 
  wire  _GEN_121; 
  wire  _GEN_131; 
  wire  _GEN_141; 
  wire  _GEN_153; 
  wire  _GEN_165; 
  wire  _GEN_171; 
  wire  _GEN_177; 
  wire  _GEN_183; 
  wire  _GEN_195; 
  wire  _GEN_205; 
  wire  _GEN_219; 
  wire  _GEN_231; 
  wire  _GEN_241; 
  wire  _GEN_249; 
  dual_plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0)) plusarg_reader ( 
    .out(plusarg_reader_out)
  );
  assign _T_7 = io_in_a_bits_source[6:4]; 
  assign _T_8 = _T_7 == 3'h0; 
  assign _T_16 = _T_7 == 3'h1; 
  assign _T_24 = _T_7 == 3'h2; 
  assign _T_32 = _T_7 == 3'h3; 
  assign _T_40 = _T_7 == 3'h4; 
  assign _T_48 = _T_7 == 3'h5; 
  assign _T_56 = _T_7 == 3'h6; 
  assign _T_64 = _T_7 == 3'h7; 
  assign _T_70 = _T_8 | _T_16; 
  assign _T_71 = _T_70 | _T_24; 
  assign _T_72 = _T_71 | _T_32; 
  assign _T_73 = _T_72 | _T_40; 
  assign _T_74 = _T_73 | _T_48; 
  assign _T_75 = _T_74 | _T_56; 
  assign _T_76 = _T_75 | _T_64; 
  assign _T_78 = 13'h3f << io_in_a_bits_size; 
  assign _T_79 = _T_78[5:0]; 
  assign _T_80 = ~ _T_79; 
  assign _GEN_33 = {{23'd0}, _T_80}; 
  assign _T_81 = io_in_a_bits_address & _GEN_33; 
  assign _T_82 = _T_81 == 29'h0; 
  assign _T_84 = io_in_a_bits_size[1:0]; 
  assign _T_85 = 4'h1 << _T_84; 
  assign _T_86 = _T_85[2:0]; 
  assign _T_87 = _T_86 | 3'h1; 
  assign _T_88 = io_in_a_bits_size >= 3'h3; 
  assign _T_89 = _T_87[2]; 
  assign _T_90 = io_in_a_bits_address[2]; 
  assign _T_91 = _T_90 == 1'h0; 
  assign _T_93 = _T_89 & _T_91; 
  assign _T_94 = _T_88 | _T_93; 
  assign _T_96 = _T_89 & _T_90; 
  assign _T_97 = _T_88 | _T_96; 
  assign _T_98 = _T_87[1]; 
  assign _T_99 = io_in_a_bits_address[1]; 
  assign _T_100 = _T_99 == 1'h0; 
  assign _T_101 = _T_91 & _T_100; 
  assign _T_102 = _T_98 & _T_101; 
  assign _T_103 = _T_94 | _T_102; 
  assign _T_104 = _T_91 & _T_99; 
  assign _T_105 = _T_98 & _T_104; 
  assign _T_106 = _T_94 | _T_105; 
  assign _T_107 = _T_90 & _T_100; 
  assign _T_108 = _T_98 & _T_107; 
  assign _T_109 = _T_97 | _T_108; 
  assign _T_110 = _T_90 & _T_99; 
  assign _T_111 = _T_98 & _T_110; 
  assign _T_112 = _T_97 | _T_111; 
  assign _T_113 = _T_87[0]; 
  assign _T_114 = io_in_a_bits_address[0]; 
  assign _T_115 = _T_114 == 1'h0; 
  assign _T_116 = _T_101 & _T_115; 
  assign _T_117 = _T_113 & _T_116; 
  assign _T_118 = _T_103 | _T_117; 
  assign _T_119 = _T_101 & _T_114; 
  assign _T_120 = _T_113 & _T_119; 
  assign _T_121 = _T_103 | _T_120; 
  assign _T_122 = _T_104 & _T_115; 
  assign _T_123 = _T_113 & _T_122; 
  assign _T_124 = _T_106 | _T_123; 
  assign _T_125 = _T_104 & _T_114; 
  assign _T_126 = _T_113 & _T_125; 
  assign _T_127 = _T_106 | _T_126; 
  assign _T_128 = _T_107 & _T_115; 
  assign _T_129 = _T_113 & _T_128; 
  assign _T_130 = _T_109 | _T_129; 
  assign _T_131 = _T_107 & _T_114; 
  assign _T_132 = _T_113 & _T_131; 
  assign _T_133 = _T_109 | _T_132; 
  assign _T_134 = _T_110 & _T_115; 
  assign _T_135 = _T_113 & _T_134; 
  assign _T_136 = _T_112 | _T_135; 
  assign _T_137 = _T_110 & _T_114; 
  assign _T_138 = _T_113 & _T_137; 
  assign _T_139 = _T_112 | _T_138; 
  assign _T_146 = {_T_139,_T_136,_T_133,_T_130,_T_127,_T_124,_T_121,_T_118}; 
  assign _T_277 = io_in_a_bits_opcode == 3'h6; 
  assign _T_279 = io_in_a_bits_size <= 3'h6; 
  assign _T_282 = io_in_a_bits_address ^ 29'h10000000; 
  assign _T_283 = {1'b0,$signed(_T_282)}; 
  assign _T_284 = $signed(_T_283) & $signed(-30'sh10000000); 
  assign _T_285 = $signed(_T_284); 
  assign _T_286 = $signed(_T_285) == $signed(30'sh0); 
  assign _T_287 = _T_279 & _T_286; 
  assign _T_290 = _T_287 | reset; 
  assign _T_291 = _T_290 == 1'h0; 
  assign _T_360 = _T_8 ? _T_279 : 1'h0; 
  assign _T_377 = _T_360 | reset; 
  assign _T_378 = _T_377 == 1'h0; 
  assign _T_380 = _T_76 | reset; 
  assign _T_381 = _T_380 == 1'h0; 
  assign _T_384 = _T_88 | reset; 
  assign _T_385 = _T_384 == 1'h0; 
  assign _T_387 = _T_82 | reset; 
  assign _T_388 = _T_387 == 1'h0; 
  assign _T_389 = io_in_a_bits_param <= 3'h2; 
  assign _T_391 = _T_389 | reset; 
  assign _T_392 = _T_391 == 1'h0; 
  assign _T_393 = ~ io_in_a_bits_mask; 
  assign _T_394 = _T_393 == 8'h0; 
  assign _T_396 = _T_394 | reset; 
  assign _T_397 = _T_396 == 1'h0; 
  assign _T_398 = io_in_a_bits_corrupt == 1'h0; 
  assign _T_400 = _T_398 | reset; 
  assign _T_401 = _T_400 == 1'h0; 
  assign _T_402 = io_in_a_bits_opcode == 3'h7; 
  assign _T_518 = io_in_a_bits_param != 3'h0; 
  assign _T_520 = _T_518 | reset; 
  assign _T_521 = _T_520 == 1'h0; 
  assign _T_531 = io_in_a_bits_opcode == 3'h4; 
  assign _T_552 = io_in_a_bits_param == 3'h0; 
  assign _T_554 = _T_552 | reset; 
  assign _T_555 = _T_554 == 1'h0; 
  assign _T_556 = io_in_a_bits_mask == _T_146; 
  assign _T_558 = _T_556 | reset; 
  assign _T_559 = _T_558 == 1'h0; 
  assign _T_564 = io_in_a_bits_opcode == 3'h0; 
  assign _T_593 = io_in_a_bits_opcode == 3'h1; 
  assign _T_618 = ~ _T_146; 
  assign _T_619 = io_in_a_bits_mask & _T_618; 
  assign _T_620 = _T_619 == 8'h0; 
  assign _T_622 = _T_620 | reset; 
  assign _T_623 = _T_622 == 1'h0; 
  assign _T_624 = io_in_a_bits_opcode == 3'h2; 
  assign _T_645 = io_in_a_bits_param <= 3'h4; 
  assign _T_647 = _T_645 | reset; 
  assign _T_648 = _T_647 == 1'h0; 
  assign _T_653 = io_in_a_bits_opcode == 3'h3; 
  assign _T_674 = io_in_a_bits_param <= 3'h3; 
  assign _T_676 = _T_674 | reset; 
  assign _T_677 = _T_676 == 1'h0; 
  assign _T_682 = io_in_a_bits_opcode == 3'h5; 
  assign _T_711 = io_in_d_bits_opcode <= 3'h6; 
  assign _T_713 = _T_711 | reset; 
  assign _T_714 = _T_713 == 1'h0; 
  assign _T_717 = io_in_d_bits_source[6:4]; 
  assign _T_718 = _T_717 == 3'h0; 
  assign _T_726 = _T_717 == 3'h1; 
  assign _T_734 = _T_717 == 3'h2; 
  assign _T_742 = _T_717 == 3'h3; 
  assign _T_750 = _T_717 == 3'h4; 
  assign _T_758 = _T_717 == 3'h5; 
  assign _T_766 = _T_717 == 3'h6; 
  assign _T_774 = _T_717 == 3'h7; 
  assign _T_780 = _T_718 | _T_726; 
  assign _T_781 = _T_780 | _T_734; 
  assign _T_782 = _T_781 | _T_742; 
  assign _T_783 = _T_782 | _T_750; 
  assign _T_784 = _T_783 | _T_758; 
  assign _T_785 = _T_784 | _T_766; 
  assign _T_786 = _T_785 | _T_774; 
  assign _T_787 = io_in_d_bits_sink < 1'h1; 
  assign _T_788 = io_in_d_bits_opcode == 3'h6; 
  assign _T_790 = _T_786 | reset; 
  assign _T_791 = _T_790 == 1'h0; 
  assign _T_792 = io_in_d_bits_size >= 3'h3; 
  assign _T_794 = _T_792 | reset; 
  assign _T_795 = _T_794 == 1'h0; 
  assign _T_796 = io_in_d_bits_param == 2'h0; 
  assign _T_798 = _T_796 | reset; 
  assign _T_799 = _T_798 == 1'h0; 
  assign _T_800 = io_in_d_bits_corrupt == 1'h0; 
  assign _T_802 = _T_800 | reset; 
  assign _T_803 = _T_802 == 1'h0; 
  assign _T_804 = io_in_d_bits_denied == 1'h0; 
  assign _T_806 = _T_804 | reset; 
  assign _T_807 = _T_806 == 1'h0; 
  assign _T_808 = io_in_d_bits_opcode == 3'h4; 
  assign _T_813 = _T_787 | reset; 
  assign _T_814 = _T_813 == 1'h0; 
  assign _T_819 = io_in_d_bits_param <= 2'h2; 
  assign _T_821 = _T_819 | reset; 
  assign _T_822 = _T_821 == 1'h0; 
  assign _T_823 = io_in_d_bits_param != 2'h2; 
  assign _T_825 = _T_823 | reset; 
  assign _T_826 = _T_825 == 1'h0; 
  assign _T_836 = io_in_d_bits_opcode == 3'h5; 
  assign _T_856 = _T_804 | io_in_d_bits_corrupt; 
  assign _T_858 = _T_856 | reset; 
  assign _T_859 = _T_858 == 1'h0; 
  assign _T_865 = io_in_d_bits_opcode == 3'h0; 
  assign _T_882 = io_in_d_bits_opcode == 3'h1; 
  assign _T_900 = io_in_d_bits_opcode == 3'h2; 
  assign _T_1456 = io_in_c_bits_source[6:4]; 
  assign _T_1457 = _T_1456 == 3'h0; 
  assign _T_1465 = _T_1456 == 3'h1; 
  assign _T_1473 = _T_1456 == 3'h2; 
  assign _T_1481 = _T_1456 == 3'h3; 
  assign _T_1489 = _T_1456 == 3'h4; 
  assign _T_1497 = _T_1456 == 3'h5; 
  assign _T_1505 = _T_1456 == 3'h6; 
  assign _T_1513 = _T_1456 == 3'h7; 
  assign _T_1519 = _T_1457 | _T_1465; 
  assign _T_1520 = _T_1519 | _T_1473; 
  assign _T_1521 = _T_1520 | _T_1481; 
  assign _T_1522 = _T_1521 | _T_1489; 
  assign _T_1523 = _T_1522 | _T_1497; 
  assign _T_1524 = _T_1523 | _T_1505; 
  assign _T_1525 = _T_1524 | _T_1513; 
  assign _T_1527 = 13'h3f << io_in_c_bits_size; 
  assign _T_1528 = _T_1527[5:0]; 
  assign _T_1529 = ~ _T_1528; 
  assign _GEN_34 = {{23'd0}, _T_1529}; 
  assign _T_1530 = io_in_c_bits_address & _GEN_34; 
  assign _T_1531 = _T_1530 == 29'h0; 
  assign _T_1532 = io_in_c_bits_address ^ 29'h10000000; 
  assign _T_1533 = {1'b0,$signed(_T_1532)}; 
  assign _T_1534 = $signed(_T_1533) & $signed(-30'sh10000000); 
  assign _T_1535 = $signed(_T_1534); 
  assign _T_1536 = $signed(_T_1535) == $signed(30'sh0); 
  assign _T_1668 = io_in_c_bits_opcode == 3'h4; 
  assign _T_1670 = _T_1536 | reset; 
  assign _T_1671 = _T_1670 == 1'h0; 
  assign _T_1673 = _T_1525 | reset; 
  assign _T_1674 = _T_1673 == 1'h0; 
  assign _T_1675 = io_in_c_bits_size >= 3'h3; 
  assign _T_1677 = _T_1675 | reset; 
  assign _T_1678 = _T_1677 == 1'h0; 
  assign _T_1680 = _T_1531 | reset; 
  assign _T_1681 = _T_1680 == 1'h0; 
  assign _T_1682 = io_in_c_bits_param <= 3'h5; 
  assign _T_1684 = _T_1682 | reset; 
  assign _T_1685 = _T_1684 == 1'h0; 
  assign _T_1686 = io_in_c_bits_corrupt == 1'h0; 
  assign _T_1688 = _T_1686 | reset; 
  assign _T_1689 = _T_1688 == 1'h0; 
  assign _T_1690 = io_in_c_bits_opcode == 3'h5; 
  assign _T_1708 = io_in_c_bits_opcode == 3'h6; 
  assign _T_1710 = io_in_c_bits_size <= 3'h6; 
  assign _T_1718 = _T_1710 & _T_1536; 
  assign _T_1721 = _T_1718 | reset; 
  assign _T_1722 = _T_1721 == 1'h0; 
  assign _T_1791 = _T_1457 ? _T_1710 : 1'h0; 
  assign _T_1808 = _T_1791 | reset; 
  assign _T_1809 = _T_1808 == 1'h0; 
  assign _T_1820 = io_in_c_bits_param <= 3'h2; 
  assign _T_1822 = _T_1820 | reset; 
  assign _T_1823 = _T_1822 == 1'h0; 
  assign _T_1828 = io_in_c_bits_opcode == 3'h7; 
  assign _T_1944 = io_in_c_bits_opcode == 3'h0; 
  assign _T_1954 = io_in_c_bits_param == 3'h0; 
  assign _T_1956 = _T_1954 | reset; 
  assign _T_1957 = _T_1956 == 1'h0; 
  assign _T_1962 = io_in_c_bits_opcode == 3'h1; 
  assign _T_1976 = io_in_c_bits_opcode == 3'h2; 
  assign _T_1998 = io_in_a_ready & io_in_a_valid; 
  assign _T_2003 = _T_80[5:3]; 
  assign _T_2004 = io_in_a_bits_opcode[2]; 
  assign _T_2005 = _T_2004 == 1'h0; 
  assign _T_2009 = _T_2007 - 3'h1; 
  assign _T_2010 = _T_2007 == 3'h0; 
  assign _T_2023 = _T_2010 == 1'h0; 
  assign _T_2024 = io_in_a_valid & _T_2023; 
  assign _T_2025 = io_in_a_bits_opcode == _T_2018; 
  assign _T_2027 = _T_2025 | reset; 
  assign _T_2028 = _T_2027 == 1'h0; 
  assign _T_2029 = io_in_a_bits_param == _T_2019; 
  assign _T_2031 = _T_2029 | reset; 
  assign _T_2032 = _T_2031 == 1'h0; 
  assign _T_2033 = io_in_a_bits_size == _T_2020; 
  assign _T_2035 = _T_2033 | reset; 
  assign _T_2036 = _T_2035 == 1'h0; 
  assign _T_2037 = io_in_a_bits_source == _T_2021; 
  assign _T_2039 = _T_2037 | reset; 
  assign _T_2040 = _T_2039 == 1'h0; 
  assign _T_2041 = io_in_a_bits_address == _T_2022; 
  assign _T_2043 = _T_2041 | reset; 
  assign _T_2044 = _T_2043 == 1'h0; 
  assign _T_2046 = _T_1998 & _T_2010; 
  assign _T_2047 = io_in_d_ready & io_in_d_valid; 
  assign _T_2049 = 13'h3f << io_in_d_bits_size; 
  assign _T_2050 = _T_2049[5:0]; 
  assign _T_2051 = ~ _T_2050; 
  assign _T_2052 = _T_2051[5:3]; 
  assign _T_2053 = io_in_d_bits_opcode[0]; 
  assign _T_2057 = _T_2055 - 3'h1; 
  assign _T_2058 = _T_2055 == 3'h0; 
  assign _T_2072 = _T_2058 == 1'h0; 
  assign _T_2073 = io_in_d_valid & _T_2072; 
  assign _T_2074 = io_in_d_bits_opcode == _T_2066; 
  assign _T_2076 = _T_2074 | reset; 
  assign _T_2077 = _T_2076 == 1'h0; 
  assign _T_2078 = io_in_d_bits_param == _T_2067; 
  assign _T_2080 = _T_2078 | reset; 
  assign _T_2081 = _T_2080 == 1'h0; 
  assign _T_2082 = io_in_d_bits_size == _T_2068; 
  assign _T_2084 = _T_2082 | reset; 
  assign _T_2085 = _T_2084 == 1'h0; 
  assign _T_2086 = io_in_d_bits_source == _T_2069; 
  assign _T_2088 = _T_2086 | reset; 
  assign _T_2089 = _T_2088 == 1'h0; 
  assign _T_2090 = io_in_d_bits_sink == _T_2070; 
  assign _T_2092 = _T_2090 | reset; 
  assign _T_2093 = _T_2092 == 1'h0; 
  assign _T_2094 = io_in_d_bits_denied == _T_2071; 
  assign _T_2096 = _T_2094 | reset; 
  assign _T_2097 = _T_2096 == 1'h0; 
  assign _T_2099 = _T_2047 & _T_2058; 
  assign _T_2149 = io_in_c_ready & io_in_c_valid; 
  assign _T_2154 = _T_1529[5:3]; 
  assign _T_2155 = io_in_c_bits_opcode[0]; 
  assign _T_2159 = _T_2157 - 3'h1; 
  assign _T_2160 = _T_2157 == 3'h0; 
  assign _T_2173 = _T_2160 == 1'h0; 
  assign _T_2174 = io_in_c_valid & _T_2173; 
  assign _T_2175 = io_in_c_bits_opcode == _T_2168; 
  assign _T_2177 = _T_2175 | reset; 
  assign _T_2178 = _T_2177 == 1'h0; 
  assign _T_2179 = io_in_c_bits_param == _T_2169; 
  assign _T_2181 = _T_2179 | reset; 
  assign _T_2182 = _T_2181 == 1'h0; 
  assign _T_2183 = io_in_c_bits_size == _T_2170; 
  assign _T_2185 = _T_2183 | reset; 
  assign _T_2186 = _T_2185 == 1'h0; 
  assign _T_2187 = io_in_c_bits_source == _T_2171; 
  assign _T_2189 = _T_2187 | reset; 
  assign _T_2190 = _T_2189 == 1'h0; 
  assign _T_2191 = io_in_c_bits_address == _T_2172; 
  assign _T_2193 = _T_2191 | reset; 
  assign _T_2194 = _T_2193 == 1'h0; 
  assign _T_2196 = _T_2149 & _T_2160; 
  assign _T_2209 = _T_2207 - 3'h1; 
  assign _T_2210 = _T_2207 == 3'h0; 
  assign _T_2228 = _T_2226 - 3'h1; 
  assign _T_2229 = _T_2226 == 3'h0; 
  assign _T_2239 = _T_1998 & _T_2210; 
  assign _T_2241 = 128'h1 << io_in_a_bits_source; 
  assign _T_2242 = _T_2197 >> io_in_a_bits_source; 
  assign _T_2243 = _T_2242[0]; 
  assign _T_2244 = _T_2243 == 1'h0; 
  assign _T_2246 = _T_2244 | reset; 
  assign _T_2247 = _T_2246 == 1'h0; 
  assign _GEN_27 = _T_2239 ? _T_2241 : 128'h0; 
  assign _T_2251 = _T_2047 & _T_2229; 
  assign _T_2253 = _T_788 == 1'h0; 
  assign _T_2254 = _T_2251 & _T_2253; 
  assign _T_2255 = 128'h1 << io_in_d_bits_source; 
  assign _T_2256 = _GEN_27 | _T_2197; 
  assign _T_2257 = _T_2256 >> io_in_d_bits_source; 
  assign _T_2258 = _T_2257[0]; 
  assign _T_2260 = _T_2258 | reset; 
  assign _T_2261 = _T_2260 == 1'h0; 
  assign _GEN_28 = _T_2254 ? _T_2255 : 128'h0; 
  assign _T_2262 = _GEN_27 != _GEN_28; 
  assign _T_2263 = _GEN_27 != 128'h0; 
  assign _T_2264 = _T_2263 == 1'h0; 
  assign _T_2265 = _T_2262 | _T_2264; 
  assign _T_2267 = _T_2265 | reset; 
  assign _T_2268 = _T_2267 == 1'h0; 
  assign _T_2269 = _T_2197 | _GEN_27; 
  assign _T_2270 = ~ _GEN_28; 
  assign _T_2271 = _T_2269 & _T_2270; 
  assign _T_2273 = _T_2197 != 128'h0; 
  assign _T_2274 = _T_2273 == 1'h0; 
  assign _T_2275 = plusarg_reader_out == 32'h0; 
  assign _T_2276 = _T_2274 | _T_2275; 
  assign _T_2277 = _T_2272 < plusarg_reader_out; 
  assign _T_2278 = _T_2276 | _T_2277; 
  assign _T_2280 = _T_2278 | reset; 
  assign _T_2281 = _T_2280 == 1'h0; 
  assign _T_2283 = _T_2272 + 32'h1; 
  assign _T_2286 = _T_1998 | _T_2047; 
  assign _T_2298 = _T_2296 - 3'h1; 
  assign _T_2299 = _T_2296 == 3'h0; 
  assign _T_2309 = _T_2047 & _T_2299; 
  assign _T_2310 = io_in_d_bits_opcode[2]; 
  assign _T_2311 = io_in_d_bits_opcode[1]; 
  assign _T_2312 = _T_2311 == 1'h0; 
  assign _T_2313 = _T_2310 & _T_2312; 
  assign _T_2314 = _T_2309 & _T_2313; 
  assign _T_2315 = 2'h1 << io_in_d_bits_sink; 
  assign _T_2316 = _T_2287 >> io_in_d_bits_sink; 
  assign _T_2318 = _T_2316 == 1'h0; 
  assign _T_2320 = _T_2318 | reset; 
  assign _T_2321 = _T_2320 == 1'h0; 
  assign _GEN_31 = _T_2314 ? _T_2315 : 2'h0; 
  assign _T_2307 = _GEN_31[0]; 
  assign _T_2327 = _T_2307 | _T_2287; 
  assign _T_2331 = _T_2327 | reset; 
  assign _T_2332 = _T_2331 == 1'h0; 
  assign _GEN_32 = io_in_e_valid ? 2'h1 : 2'h0; 
  assign _T_2333 = _T_2287 | _T_2307; 
  assign _T_2322 = _GEN_32[0]; 
  assign _T_2334 = ~ _T_2322; 
  assign _T_2335 = _T_2333 & _T_2334; 
  assign _GEN_35 = io_in_a_valid & _T_277; 
  assign _GEN_51 = io_in_a_valid & _T_402; 
  assign _GEN_69 = io_in_a_valid & _T_531; 
  assign _GEN_81 = io_in_a_valid & _T_564; 
  assign _GEN_91 = io_in_a_valid & _T_593; 
  assign _GEN_101 = io_in_a_valid & _T_624; 
  assign _GEN_111 = io_in_a_valid & _T_653; 
  assign _GEN_121 = io_in_a_valid & _T_682; 
  assign _GEN_131 = io_in_d_valid & _T_788; 
  assign _GEN_141 = io_in_d_valid & _T_808; 
  assign _GEN_153 = io_in_d_valid & _T_836; 
  assign _GEN_165 = io_in_d_valid & _T_865; 
  assign _GEN_171 = io_in_d_valid & _T_882; 
  assign _GEN_177 = io_in_d_valid & _T_900; 
  assign _GEN_183 = io_in_c_valid & _T_1668; 
  assign _GEN_195 = io_in_c_valid & _T_1690; 
  assign _GEN_205 = io_in_c_valid & _T_1708; 
  assign _GEN_219 = io_in_c_valid & _T_1828; 
  assign _GEN_231 = io_in_c_valid & _T_1944; 
  assign _GEN_241 = io_in_c_valid & _T_1962; 
  assign _GEN_249 = io_in_c_valid & _T_1976; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2007 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_2018 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2019 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_2020 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_2021 = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_2022 = _RAND_5[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_2055 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_2066 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_2067 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_2068 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_2069 = _RAND_10[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_2070 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_2071 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_2157 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_2168 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_2169 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_2170 = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_2171 = _RAND_17[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_2172 = _RAND_18[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {4{`RANDOM}};
  _T_2197 = _RAND_19[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_2207 = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_2226 = _RAND_21[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_2272 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_2287 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_2296 = _RAND_24[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_2007 <= 3'h0;
    end else begin
      if (_T_1998) begin
        if (_T_2010) begin
          if (_T_2005) begin
            _T_2007 <= _T_2003;
          end else begin
            _T_2007 <= 3'h0;
          end
        end else begin
          _T_2007 <= _T_2009;
        end
      end
    end
    if (_T_2046) begin
      _T_2018 <= io_in_a_bits_opcode;
    end
    if (_T_2046) begin
      _T_2019 <= io_in_a_bits_param;
    end
    if (_T_2046) begin
      _T_2020 <= io_in_a_bits_size;
    end
    if (_T_2046) begin
      _T_2021 <= io_in_a_bits_source;
    end
    if (_T_2046) begin
      _T_2022 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_2055 <= 3'h0;
    end else begin
      if (_T_2047) begin
        if (_T_2058) begin
          if (_T_2053) begin
            _T_2055 <= _T_2052;
          end else begin
            _T_2055 <= 3'h0;
          end
        end else begin
          _T_2055 <= _T_2057;
        end
      end
    end
    if (_T_2099) begin
      _T_2066 <= io_in_d_bits_opcode;
    end
    if (_T_2099) begin
      _T_2067 <= io_in_d_bits_param;
    end
    if (_T_2099) begin
      _T_2068 <= io_in_d_bits_size;
    end
    if (_T_2099) begin
      _T_2069 <= io_in_d_bits_source;
    end
    if (_T_2099) begin
      _T_2070 <= io_in_d_bits_sink;
    end
    if (_T_2099) begin
      _T_2071 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_2157 <= 3'h0;
    end else begin
      if (_T_2149) begin
        if (_T_2160) begin
          if (_T_2155) begin
            _T_2157 <= _T_2154;
          end else begin
            _T_2157 <= 3'h0;
          end
        end else begin
          _T_2157 <= _T_2159;
        end
      end
    end
    if (_T_2196) begin
      _T_2168 <= io_in_c_bits_opcode;
    end
    if (_T_2196) begin
      _T_2169 <= io_in_c_bits_param;
    end
    if (_T_2196) begin
      _T_2170 <= io_in_c_bits_size;
    end
    if (_T_2196) begin
      _T_2171 <= io_in_c_bits_source;
    end
    if (_T_2196) begin
      _T_2172 <= io_in_c_bits_address;
    end
    if (reset) begin
      _T_2197 <= 128'h0;
    end else begin
      _T_2197 <= _T_2271;
    end
    if (reset) begin
      _T_2207 <= 3'h0;
    end else begin
      if (_T_1998) begin
        if (_T_2210) begin
          if (_T_2005) begin
            _T_2207 <= _T_2003;
          end else begin
            _T_2207 <= 3'h0;
          end
        end else begin
          _T_2207 <= _T_2209;
        end
      end
    end
    if (reset) begin
      _T_2226 <= 3'h0;
    end else begin
      if (_T_2047) begin
        if (_T_2229) begin
          if (_T_2053) begin
            _T_2226 <= _T_2052;
          end else begin
            _T_2226 <= 3'h0;
          end
        end else begin
          _T_2226 <= _T_2228;
        end
      end
    end
    if (reset) begin
      _T_2272 <= 32'h0;
    end else begin
      if (_T_2286) begin
        _T_2272 <= 32'h0;
      end else begin
        _T_2272 <= _T_2283;
      end
    end
    if (reset) begin
      _T_2287 <= 1'h0;
    end else begin
      _T_2287 <= _T_2335;
    end
    if (reset) begin
      _T_2296 <= 3'h0;
    end else begin
      if (_T_2047) begin
        if (_T_2299) begin
          if (_T_2053) begin
            _T_2296 <= _T_2052;
          end else begin
            _T_2296 <= 3'h0;
          end
        end else begin
          _T_2296 <= _T_2298;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel has invalid opcode (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:39 assert (TLMessages.isA(bundle.opcode), \"'A' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:46 assert (visible(edge.address(bundle), bundle.source, edge), \"'A' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_291) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_291) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_378) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_378) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_381) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_381) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_385) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_388) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_388) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_392) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_392) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_397) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_397) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_401) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:56 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_401) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_291) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_291) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_378) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_378) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_381) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_381) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_385) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_388) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_388) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_392) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_392) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_521) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_521) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_397) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_397) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_401) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:68 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_401) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_291) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & _T_291) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_381) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & _T_381) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_388) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & _T_388) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_555) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & _T_555) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_559) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & _T_559) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_401) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:77 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & _T_401) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_81 & _T_291) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_81 & _T_291) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_81 & _T_381) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_81 & _T_381) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_81 & _T_388) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_81 & _T_388) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_81 & _T_555) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_81 & _T_555) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_81 & _T_559) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_81 & _T_559) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_291) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_291) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_381) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_381) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_388) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_388) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_555) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_555) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_623) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_623) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_291) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_291) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_381) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_381) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_388) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_388) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_648) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_648) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_559) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_559) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & _T_291) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & _T_291) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & _T_381) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & _T_381) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & _T_388) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & _T_388) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & _T_677) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & _T_677) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & _T_559) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & _T_559) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_291) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_291) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_381) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_381) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_388) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_388) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_559) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_559) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_401) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:117 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_401) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_714) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_714) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_791) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_791) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_795) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_795) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_799) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_799) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_803) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_803) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_807) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_807) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_791) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_791) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_814) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:285 assert (sink_ok, \"'D' channel Grant carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_814) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_795) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_795) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_822) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_822) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_826) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_826) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_803) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_803) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is denied (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:290 assert (deny_put_ok || !bundle.denied, \"'D' channel Grant is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_791) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_791) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_814) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:295 assert (sink_ok, \"'D' channel GrantData carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_814) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_795) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_795) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_822) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_822) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_826) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_826) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_859) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_859) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:300 assert (deny_get_ok || !bundle.denied, \"'D' channel GrantData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & _T_791) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & _T_791) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & _T_799) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & _T_799) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & _T_803) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & _T_803) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is denied (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:308 assert (deny_put_ok || !bundle.denied, \"'D' channel AccessAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_791) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_791) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_799) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_799) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_859) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_859) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:316 assert (deny_get_ok || !bundle.denied, \"'D' channel AccessAckData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_177 & _T_791) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_177 & _T_791) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_177 & _T_799) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_177 & _T_799) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_177 & _T_803) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_177 & _T_803) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is denied (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:324 assert (deny_put_ok || !bundle.denied, \"'D' channel HintAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel has invalid opcode (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:122 assert (TLMessages.isB(bundle.opcode), \"'B' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:124 assert (visible(edge.address(bundle), bundle.source, edge), \"'B' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Probe type unsupported by client (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:133 assert (edge.client.supportsProbe(bundle.source, bundle.size), \"'B' channel carries Probe type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:134 assert (address_ok, \"'B' channel Probe carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries source that is not first source (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:135 assert (legal_source, \"'B' channel Probe carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:136 assert (is_aligned, \"'B' channel Probe address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:137 assert (TLPermissions.isCap(bundle.param), \"'B' channel Probe carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe contains invalid mask (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:138 assert (bundle.mask === mask, \"'B' channel Probe contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe is corrupt (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:139 assert (!bundle.corrupt, \"'B' channel Probe is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Get type unsupported by client (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:143 assert (edge.client.supportsGet(bundle.source, bundle.size), \"'B' channel carries Get type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries unmanaged address (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:144 assert (address_ok, \"'B' channel Get carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries source that is not first source (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:145 assert (legal_source, \"'B' channel Get carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:146 assert (is_aligned, \"'B' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries invalid param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:147 assert (bundle.param === UInt(0), \"'B' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get contains invalid mask (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:148 assert (bundle.mask === mask, \"'B' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get is corrupt (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:149 assert (!bundle.corrupt, \"'B' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutFull type unsupported by client (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:153 assert (edge.client.supportsPutFull(bundle.source, bundle.size), \"'B' channel carries PutFull type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries unmanaged address (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:154 assert (address_ok, \"'B' channel PutFull carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries source that is not first source (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:155 assert (legal_source, \"'B' channel PutFull carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:156 assert (is_aligned, \"'B' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries invalid param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:157 assert (bundle.param === UInt(0), \"'B' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull contains invalid mask (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:158 assert (bundle.mask === mask, \"'B' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutPartial type unsupported by client (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:162 assert (edge.client.supportsPutPartial(bundle.source, bundle.size), \"'B' channel carries PutPartial type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:163 assert (address_ok, \"'B' channel PutPartial carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:164 assert (legal_source, \"'B' channel PutPartial carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:165 assert (is_aligned, \"'B' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries invalid param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:166 assert (bundle.param === UInt(0), \"'B' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial contains invalid mask (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:167 assert ((bundle.mask & ~mask) === UInt(0), \"'B' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Arithmetic type unsupported by client (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:171 assert (edge.client.supportsArithmetic(bundle.source, bundle.size), \"'B' channel carries Arithmetic type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:172 assert (address_ok, \"'B' channel Arithmetic carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:173 assert (legal_source, \"'B' channel Arithmetic carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:174 assert (is_aligned, \"'B' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries invalid opcode param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:175 assert (TLAtomics.isArithmetic(bundle.param), \"'B' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:176 assert (bundle.mask === mask, \"'B' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Logical type unsupported by client (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:180 assert (edge.client.supportsLogical(bundle.source, bundle.size), \"'B' channel carries Logical type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries unmanaged address (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:181 assert (address_ok, \"'B' channel Logical carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries source that is not first source (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:182 assert (legal_source, \"'B' channel Logical carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:183 assert (is_aligned, \"'B' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries invalid opcode param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:184 assert (TLAtomics.isLogical(bundle.param), \"'B' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical contains invalid mask (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:185 assert (bundle.mask === mask, \"'B' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Hint type unsupported by client (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:189 assert (edge.client.supportsHint(bundle.source, bundle.size), \"'B' channel carries Hint type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries unmanaged address (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:190 assert (address_ok, \"'B' channel Hint carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries source that is not first source (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:191 assert (legal_source, \"'B' channel Hint carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:192 assert (is_aligned, \"'B' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint contains invalid mask (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:193 assert (bundle.mask === mask, \"'B' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint is corrupt (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:194 assert (!bundle.corrupt, \"'B' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel has invalid opcode (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:199 assert (TLMessages.isC(bundle.opcode), \"'C' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:205 assert (visible(edge.address(bundle), bundle.source, edge), \"'C' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_1671) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:208 assert (address_ok, \"'C' channel ProbeAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_1671) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_1674) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:209 assert (source_ok, \"'C' channel ProbeAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_1674) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_1678) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:210 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_1678) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_1681) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:211 assert (is_aligned, \"'C' channel ProbeAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_1681) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_1685) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:212 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAck carries invalid report param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_1685) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_1689) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck is corrupt (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:213 assert (!bundle.corrupt, \"'C' channel ProbeAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_1689) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1671) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:217 assert (address_ok, \"'C' channel ProbeAckData carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1671) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1674) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:218 assert (source_ok, \"'C' channel ProbeAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1674) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1678) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:219 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAckData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1678) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1681) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:220 assert (is_aligned, \"'C' channel ProbeAckData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1681) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1685) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:221 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAckData carries invalid report param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1685) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1722) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:225 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries Release type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1722) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1809) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:226 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1809) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1674) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:227 assert (source_ok, \"'C' channel Release carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1674) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1678) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:228 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel Release smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1678) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1681) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:229 assert (is_aligned, \"'C' channel Release address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1681) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1823) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid shrink param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:230 assert (TLPermissions.isShrink(bundle.param), \"'C' channel Release carries invalid shrink param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1823) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1689) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release is corrupt (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:231 assert (!bundle.corrupt, \"'C' channel Release is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1689) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1722) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:235 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries ReleaseData type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1722) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1809) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:236 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1809) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1674) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:237 assert (source_ok, \"'C' channel ReleaseData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1674) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1678) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:238 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ReleaseData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1678) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1681) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:239 assert (is_aligned, \"'C' channel ReleaseData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1681) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1823) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid shrink param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:240 assert (TLPermissions.isShrink(bundle.param), \"'C' channel ReleaseData carries invalid shrink param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1823) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1671) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:244 assert (address_ok, \"'C' channel AccessAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1671) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1674) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:245 assert (source_ok, \"'C' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1674) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1681) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:246 assert (is_aligned, \"'C' channel AccessAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1681) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1957) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:247 assert (bundle.param === UInt(0), \"'C' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1957) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1689) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck is corrupt (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:248 assert (!bundle.corrupt, \"'C' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1689) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1671) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:252 assert (address_ok, \"'C' channel AccessAckData carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1671) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1674) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:253 assert (source_ok, \"'C' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1674) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1681) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:254 assert (is_aligned, \"'C' channel AccessAckData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1681) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1957) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:255 assert (bundle.param === UInt(0), \"'C' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1957) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_249 & _T_1671) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:259 assert (address_ok, \"'C' channel HintAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_249 & _T_1671) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_249 & _T_1674) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:260 assert (source_ok, \"'C' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_249 & _T_1674) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_249 & _T_1681) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:261 assert (is_aligned, \"'C' channel HintAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_249 & _T_1681) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_249 & _T_1957) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:262 assert (bundle.param === UInt(0), \"'C' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_249 & _T_1957) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_249 & _T_1689) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck is corrupt (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:263 assert (!bundle.corrupt, \"'C' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_249 & _T_1689) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channels carries invalid sink ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:330 assert (sink_ok, \"'E' channels carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2024 & _T_2028) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2024 & _T_2028) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2024 & _T_2032) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2024 & _T_2032) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2024 & _T_2036) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2024 & _T_2036) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2024 & _T_2040) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2024 & _T_2040) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2024 & _T_2044) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2024 & _T_2044) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2073 & _T_2077) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2073 & _T_2077) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2073 & _T_2081) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2073 & _T_2081) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2073 & _T_2085) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2073 & _T_2085) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2073 & _T_2089) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2073 & _T_2089) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2073 & _T_2093) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2073 & _T_2093) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2073 & _T_2097) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2073 & _T_2097) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:378 assert (b.bits.opcode === opcode, \"'B' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:379 assert (b.bits.param  === param,  \"'B' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel size changed within multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:380 assert (b.bits.size   === size,   \"'B' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel source changed within multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:381 assert (b.bits.source === source, \"'B' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:382 assert (b.bits.address=== address,\"'B' channel addresss changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2174 & _T_2178) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:401 assert (c.bits.opcode === opcode, \"'C' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2174 & _T_2178) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2174 & _T_2182) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:402 assert (c.bits.param  === param,  \"'C' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2174 & _T_2182) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2174 & _T_2186) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:403 assert (c.bits.size   === size,   \"'C' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2174 & _T_2186) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2174 & _T_2190) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:404 assert (c.bits.source === source, \"'C' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2174 & _T_2190) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2174 & _T_2194) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:405 assert (c.bits.address=== address,\"'C' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2174 & _T_2194) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2239 & _T_2247) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2239 & _T_2247) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2254 & _T_2261) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2254 & _T_2261) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2268) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2268) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2281) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:479 assert (!inflight.orR || limit === UInt(0) || watchdog < limit, \"TileLink timeout expired\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2281) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2314 & _T_2321) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:494 assert(!inflight(bundle.d.bits.sink), \"'D' channel re-used a sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2314 & _T_2321) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_e_valid & _T_2332) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at ChiplinkTest.scala:363:32)\n    at Monitor.scala:500 assert((d_set | inflight)(bundle.e.bits.sink), \"'E' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_e_valid & _T_2332) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLMonitor_1( 
  input         clock, 
  input         reset, 
  input         io_in_a_ready, 
  input         io_in_a_valid, 
  input  [2:0]  io_in_a_bits_opcode, 
  input  [2:0]  io_in_a_bits_param, 
  input  [2:0]  io_in_a_bits_size, 
  input  [2:0]  io_in_a_bits_source, 
  input  [31:0] io_in_a_bits_address, 
  input  [3:0]  io_in_a_bits_mask, 
  input         io_in_a_bits_corrupt, 
  input         io_in_d_ready, 
  input         io_in_d_valid, 
  input  [2:0]  io_in_d_bits_opcode, 
  input  [1:0]  io_in_d_bits_param, 
  input  [2:0]  io_in_d_bits_size, 
  input  [2:0]  io_in_d_bits_source, 
  input  [5:0]  io_in_d_bits_sink, 
  input         io_in_d_bits_denied, 
  input         io_in_d_bits_corrupt 
);
  wire [31:0] plusarg_reader_out; 
  wire  _T_7; 
  wire  _T_8; 
  wire  _T_22; 
  wire [12:0] _T_24; 
  wire [5:0] _T_25; 
  wire [5:0] _T_26; 
  wire [31:0] _GEN_18; 
  wire [31:0] _T_27; 
  wire  _T_28; 
  wire  _T_30; 
  wire [1:0] _T_31; 
  wire [1:0] _T_33; 
  wire  _T_34; 
  wire  _T_35; 
  wire  _T_36; 
  wire  _T_37; 
  wire  _T_39; 
  wire  _T_40; 
  wire  _T_42; 
  wire  _T_43; 
  wire  _T_44; 
  wire  _T_45; 
  wire  _T_46; 
  wire  _T_47; 
  wire  _T_48; 
  wire  _T_49; 
  wire  _T_50; 
  wire  _T_51; 
  wire  _T_52; 
  wire  _T_53; 
  wire  _T_54; 
  wire  _T_55; 
  wire  _T_56; 
  wire  _T_57; 
  wire  _T_58; 
  wire [3:0] _T_61; 
  wire  _T_96; 
  wire [31:0] _T_98; 
  wire [32:0] _T_99; 
  wire [32:0] _T_100; 
  wire [32:0] _T_101; 
  wire  _T_102; 
  wire  _T_104; 
  wire [31:0] _T_106; 
  wire [32:0] _T_107; 
  wire [32:0] _T_108; 
  wire [32:0] _T_109; 
  wire  _T_110; 
  wire  _T_111; 
  wire  _T_113; 
  wire [31:0] _T_116; 
  wire [32:0] _T_117; 
  wire [32:0] _T_118; 
  wire [32:0] _T_119; 
  wire  _T_120; 
  wire  _T_121; 
  wire  _T_124; 
  wire  _T_126; 
  wire  _T_127; 
  wire  _T_130; 
  wire  _T_132; 
  wire  _T_133; 
  wire  _T_136; 
  wire  _T_137; 
  wire  _T_139; 
  wire  _T_140; 
  wire  _T_141; 
  wire  _T_143; 
  wire  _T_144; 
  wire [3:0] _T_145; 
  wire  _T_146; 
  wire  _T_148; 
  wire  _T_149; 
  wire  _T_150; 
  wire  _T_152; 
  wire  _T_153; 
  wire  _T_154; 
  wire  _T_203; 
  wire  _T_205; 
  wire  _T_206; 
  wire  _T_216; 
  wire  _T_236; 
  wire  _T_237; 
  wire  _T_238; 
  wire  _T_241; 
  wire  _T_242; 
  wire  _T_249; 
  wire  _T_251; 
  wire  _T_252; 
  wire  _T_253; 
  wire  _T_255; 
  wire  _T_256; 
  wire  _T_261; 
  wire  _T_302; 
  wire [3:0] _T_339; 
  wire [3:0] _T_340; 
  wire  _T_341; 
  wire  _T_343; 
  wire  _T_344; 
  wire  _T_345; 
  wire  _T_347; 
  wire  _T_361; 
  wire  _T_373; 
  wire  _T_375; 
  wire  _T_376; 
  wire  _T_383; 
  wire  _T_385; 
  wire  _T_386; 
  wire  _T_391; 
  wire  _T_429; 
  wire  _T_431; 
  wire  _T_432; 
  wire  _T_437; 
  wire  _T_478; 
  wire  _T_480; 
  wire  _T_481; 
  wire  _T_484; 
  wire  _T_485; 
  wire  _T_499; 
  wire  _T_500; 
  wire  _T_501; 
  wire  _T_503; 
  wire  _T_504; 
  wire  _T_505; 
  wire  _T_507; 
  wire  _T_508; 
  wire  _T_509; 
  wire  _T_511; 
  wire  _T_512; 
  wire  _T_513; 
  wire  _T_515; 
  wire  _T_516; 
  wire  _T_517; 
  wire  _T_519; 
  wire  _T_520; 
  wire  _T_521; 
  wire  _T_526; 
  wire  _T_527; 
  wire  _T_532; 
  wire  _T_534; 
  wire  _T_535; 
  wire  _T_536; 
  wire  _T_538; 
  wire  _T_539; 
  wire  _T_549; 
  wire  _T_569; 
  wire  _T_571; 
  wire  _T_572; 
  wire  _T_578; 
  wire  _T_595; 
  wire  _T_613; 
  wire  _T_642; 
  wire [3:0] _T_647; 
  wire  _T_648; 
  wire  _T_649; 
  reg [3:0] _T_651; 
  reg [31:0] _RAND_0;
  wire [3:0] _T_653; 
  wire  _T_654; 
  reg [2:0] _T_662; 
  reg [31:0] _RAND_1;
  reg [2:0] _T_663; 
  reg [31:0] _RAND_2;
  reg [2:0] _T_664; 
  reg [31:0] _RAND_3;
  reg [2:0] _T_665; 
  reg [31:0] _RAND_4;
  reg [31:0] _T_666; 
  reg [31:0] _RAND_5;
  wire  _T_667; 
  wire  _T_668; 
  wire  _T_669; 
  wire  _T_671; 
  wire  _T_672; 
  wire  _T_673; 
  wire  _T_675; 
  wire  _T_676; 
  wire  _T_677; 
  wire  _T_679; 
  wire  _T_680; 
  wire  _T_681; 
  wire  _T_683; 
  wire  _T_684; 
  wire  _T_685; 
  wire  _T_687; 
  wire  _T_688; 
  wire  _T_690; 
  wire  _T_691; 
  wire [12:0] _T_693; 
  wire [5:0] _T_694; 
  wire [5:0] _T_695; 
  wire [3:0] _T_696; 
  wire  _T_697; 
  reg [3:0] _T_699; 
  reg [31:0] _RAND_6;
  wire [3:0] _T_701; 
  wire  _T_702; 
  reg [2:0] _T_710; 
  reg [31:0] _RAND_7;
  reg [1:0] _T_711; 
  reg [31:0] _RAND_8;
  reg [2:0] _T_712; 
  reg [31:0] _RAND_9;
  reg [2:0] _T_713; 
  reg [31:0] _RAND_10;
  reg [5:0] _T_714; 
  reg [31:0] _RAND_11;
  reg  _T_715; 
  reg [31:0] _RAND_12;
  wire  _T_716; 
  wire  _T_717; 
  wire  _T_718; 
  wire  _T_720; 
  wire  _T_721; 
  wire  _T_722; 
  wire  _T_724; 
  wire  _T_725; 
  wire  _T_726; 
  wire  _T_728; 
  wire  _T_729; 
  wire  _T_730; 
  wire  _T_732; 
  wire  _T_733; 
  wire  _T_734; 
  wire  _T_736; 
  wire  _T_737; 
  wire  _T_738; 
  wire  _T_740; 
  wire  _T_741; 
  wire  _T_743; 
  reg [7:0] _T_744; 
  reg [31:0] _RAND_13;
  reg [3:0] _T_754; 
  reg [31:0] _RAND_14;
  wire [3:0] _T_756; 
  wire  _T_757; 
  reg [3:0] _T_773; 
  reg [31:0] _RAND_15;
  wire [3:0] _T_775; 
  wire  _T_776; 
  wire  _T_786; 
  wire [7:0] _T_788; 
  wire [7:0] _T_789; 
  wire  _T_790; 
  wire  _T_791; 
  wire  _T_793; 
  wire  _T_794; 
  wire [7:0] _GEN_15; 
  wire  _T_798; 
  wire  _T_800; 
  wire  _T_801; 
  wire [7:0] _T_802; 
  wire [7:0] _T_803; 
  wire [7:0] _T_804; 
  wire  _T_805; 
  wire  _T_807; 
  wire  _T_808; 
  wire [7:0] _GEN_16; 
  wire  _T_809; 
  wire  _T_810; 
  wire  _T_811; 
  wire  _T_812; 
  wire  _T_814; 
  wire  _T_815; 
  wire [7:0] _T_816; 
  wire [7:0] _T_817; 
  wire [7:0] _T_818; 
  reg [31:0] _T_819; 
  reg [31:0] _RAND_16;
  wire  _T_820; 
  wire  _T_821; 
  wire  _T_822; 
  wire  _T_823; 
  wire  _T_824; 
  wire  _T_825; 
  wire  _T_827; 
  wire  _T_828; 
  wire [31:0] _T_830; 
  wire  _T_833; 
  wire  _GEN_19; 
  wire  _GEN_35; 
  wire  _GEN_53; 
  wire  _GEN_65; 
  wire  _GEN_75; 
  wire  _GEN_85; 
  wire  _GEN_95; 
  wire  _GEN_105; 
  wire  _GEN_115; 
  wire  _GEN_125; 
  wire  _GEN_137; 
  wire  _GEN_149; 
  wire  _GEN_155; 
  wire  _GEN_161; 
  dual_plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0)) plusarg_reader ( 
    .out(plusarg_reader_out)
  );
  assign _T_7 = io_in_a_bits_source[2:2]; 
  assign _T_8 = _T_7 == 1'h0; 
  assign _T_22 = _T_8 | _T_7; 
  assign _T_24 = 13'h3f << io_in_a_bits_size; 
  assign _T_25 = _T_24[5:0]; 
  assign _T_26 = ~ _T_25; 
  assign _GEN_18 = {{26'd0}, _T_26}; 
  assign _T_27 = io_in_a_bits_address & _GEN_18; 
  assign _T_28 = _T_27 == 32'h0; 
  assign _T_30 = io_in_a_bits_size[0]; 
  assign _T_31 = 2'h1 << _T_30; 
  assign _T_33 = _T_31 | 2'h1; 
  assign _T_34 = io_in_a_bits_size >= 3'h2; 
  assign _T_35 = _T_33[1]; 
  assign _T_36 = io_in_a_bits_address[1]; 
  assign _T_37 = _T_36 == 1'h0; 
  assign _T_39 = _T_35 & _T_37; 
  assign _T_40 = _T_34 | _T_39; 
  assign _T_42 = _T_35 & _T_36; 
  assign _T_43 = _T_34 | _T_42; 
  assign _T_44 = _T_33[0]; 
  assign _T_45 = io_in_a_bits_address[0]; 
  assign _T_46 = _T_45 == 1'h0; 
  assign _T_47 = _T_37 & _T_46; 
  assign _T_48 = _T_44 & _T_47; 
  assign _T_49 = _T_40 | _T_48; 
  assign _T_50 = _T_37 & _T_45; 
  assign _T_51 = _T_44 & _T_50; 
  assign _T_52 = _T_40 | _T_51; 
  assign _T_53 = _T_36 & _T_46; 
  assign _T_54 = _T_44 & _T_53; 
  assign _T_55 = _T_43 | _T_54; 
  assign _T_56 = _T_36 & _T_45; 
  assign _T_57 = _T_44 & _T_56; 
  assign _T_58 = _T_43 | _T_57; 
  assign _T_61 = {_T_58,_T_55,_T_52,_T_49}; 
  assign _T_96 = io_in_a_bits_opcode == 3'h6; 
  assign _T_98 = io_in_a_bits_address ^ 32'h40000000; 
  assign _T_99 = {1'b0,$signed(_T_98)}; 
  assign _T_100 = $signed(_T_99) & $signed(-33'sh20000000); 
  assign _T_101 = $signed(_T_100); 
  assign _T_102 = $signed(_T_101) == $signed(33'sh0); 
  assign _T_104 = 3'h6 == io_in_a_bits_size; 
  assign _T_106 = io_in_a_bits_address ^ 32'h80000000; 
  assign _T_107 = {1'b0,$signed(_T_106)}; 
  assign _T_108 = $signed(_T_107) & $signed(-33'sh80000000); 
  assign _T_109 = $signed(_T_108); 
  assign _T_110 = $signed(_T_109) == $signed(33'sh0); 
  assign _T_111 = _T_104 & _T_110; 
  assign _T_113 = io_in_a_bits_size <= 3'h6; 
  assign _T_116 = io_in_a_bits_address ^ 32'h10000000; 
  assign _T_117 = {1'b0,$signed(_T_116)}; 
  assign _T_118 = $signed(_T_117) & $signed(-33'sh10000000); 
  assign _T_119 = $signed(_T_118); 
  assign _T_120 = $signed(_T_119) == $signed(33'sh0); 
  assign _T_121 = _T_113 & _T_120; 
  assign _T_124 = _T_111 | _T_121; 
  assign _T_126 = _T_124 | reset; 
  assign _T_127 = _T_126 == 1'h0; 
  assign _T_130 = reset == 1'h0; 
  assign _T_132 = _T_22 | reset; 
  assign _T_133 = _T_132 == 1'h0; 
  assign _T_136 = _T_34 | reset; 
  assign _T_137 = _T_136 == 1'h0; 
  assign _T_139 = _T_28 | reset; 
  assign _T_140 = _T_139 == 1'h0; 
  assign _T_141 = io_in_a_bits_param <= 3'h2; 
  assign _T_143 = _T_141 | reset; 
  assign _T_144 = _T_143 == 1'h0; 
  assign _T_145 = ~ io_in_a_bits_mask; 
  assign _T_146 = _T_145 == 4'h0; 
  assign _T_148 = _T_146 | reset; 
  assign _T_149 = _T_148 == 1'h0; 
  assign _T_150 = io_in_a_bits_corrupt == 1'h0; 
  assign _T_152 = _T_150 | reset; 
  assign _T_153 = _T_152 == 1'h0; 
  assign _T_154 = io_in_a_bits_opcode == 3'h7; 
  assign _T_203 = io_in_a_bits_param != 3'h0; 
  assign _T_205 = _T_203 | reset; 
  assign _T_206 = _T_205 == 1'h0; 
  assign _T_216 = io_in_a_bits_opcode == 3'h4; 
  assign _T_236 = _T_102 | _T_110; 
  assign _T_237 = _T_236 | _T_120; 
  assign _T_238 = _T_113 & _T_237; 
  assign _T_241 = _T_238 | reset; 
  assign _T_242 = _T_241 == 1'h0; 
  assign _T_249 = io_in_a_bits_param == 3'h0; 
  assign _T_251 = _T_249 | reset; 
  assign _T_252 = _T_251 == 1'h0; 
  assign _T_253 = io_in_a_bits_mask == _T_61; 
  assign _T_255 = _T_253 | reset; 
  assign _T_256 = _T_255 == 1'h0; 
  assign _T_261 = io_in_a_bits_opcode == 3'h0; 
  assign _T_302 = io_in_a_bits_opcode == 3'h1; 
  assign _T_339 = ~ _T_61; 
  assign _T_340 = io_in_a_bits_mask & _T_339; 
  assign _T_341 = _T_340 == 4'h0; 
  assign _T_343 = _T_341 | reset; 
  assign _T_344 = _T_343 == 1'h0; 
  assign _T_345 = io_in_a_bits_opcode == 3'h2; 
  assign _T_347 = io_in_a_bits_size <= 3'h3; 
  assign _T_361 = _T_347 & _T_236; 
  assign _T_373 = _T_361 | _T_121; 
  assign _T_375 = _T_373 | reset; 
  assign _T_376 = _T_375 == 1'h0; 
  assign _T_383 = io_in_a_bits_param <= 3'h4; 
  assign _T_385 = _T_383 | reset; 
  assign _T_386 = _T_385 == 1'h0; 
  assign _T_391 = io_in_a_bits_opcode == 3'h3; 
  assign _T_429 = io_in_a_bits_param <= 3'h3; 
  assign _T_431 = _T_429 | reset; 
  assign _T_432 = _T_431 == 1'h0; 
  assign _T_437 = io_in_a_bits_opcode == 3'h5; 
  assign _T_478 = io_in_d_bits_opcode <= 3'h6; 
  assign _T_480 = _T_478 | reset; 
  assign _T_481 = _T_480 == 1'h0; 
  assign _T_484 = io_in_d_bits_source[2:2]; 
  assign _T_485 = _T_484 == 1'h0; 
  assign _T_499 = _T_485 | _T_484; 
  assign _T_500 = io_in_d_bits_sink < 6'h21; 
  assign _T_501 = io_in_d_bits_opcode == 3'h6; 
  assign _T_503 = _T_499 | reset; 
  assign _T_504 = _T_503 == 1'h0; 
  assign _T_505 = io_in_d_bits_size >= 3'h2; 
  assign _T_507 = _T_505 | reset; 
  assign _T_508 = _T_507 == 1'h0; 
  assign _T_509 = io_in_d_bits_param == 2'h0; 
  assign _T_511 = _T_509 | reset; 
  assign _T_512 = _T_511 == 1'h0; 
  assign _T_513 = io_in_d_bits_corrupt == 1'h0; 
  assign _T_515 = _T_513 | reset; 
  assign _T_516 = _T_515 == 1'h0; 
  assign _T_517 = io_in_d_bits_denied == 1'h0; 
  assign _T_519 = _T_517 | reset; 
  assign _T_520 = _T_519 == 1'h0; 
  assign _T_521 = io_in_d_bits_opcode == 3'h4; 
  assign _T_526 = _T_500 | reset; 
  assign _T_527 = _T_526 == 1'h0; 
  assign _T_532 = io_in_d_bits_param <= 2'h2; 
  assign _T_534 = _T_532 | reset; 
  assign _T_535 = _T_534 == 1'h0; 
  assign _T_536 = io_in_d_bits_param != 2'h2; 
  assign _T_538 = _T_536 | reset; 
  assign _T_539 = _T_538 == 1'h0; 
  assign _T_549 = io_in_d_bits_opcode == 3'h5; 
  assign _T_569 = _T_517 | io_in_d_bits_corrupt; 
  assign _T_571 = _T_569 | reset; 
  assign _T_572 = _T_571 == 1'h0; 
  assign _T_578 = io_in_d_bits_opcode == 3'h0; 
  assign _T_595 = io_in_d_bits_opcode == 3'h1; 
  assign _T_613 = io_in_d_bits_opcode == 3'h2; 
  assign _T_642 = io_in_a_ready & io_in_a_valid; 
  assign _T_647 = _T_26[5:2]; 
  assign _T_648 = io_in_a_bits_opcode[2]; 
  assign _T_649 = _T_648 == 1'h0; 
  assign _T_653 = _T_651 - 4'h1; 
  assign _T_654 = _T_651 == 4'h0; 
  assign _T_667 = _T_654 == 1'h0; 
  assign _T_668 = io_in_a_valid & _T_667; 
  assign _T_669 = io_in_a_bits_opcode == _T_662; 
  assign _T_671 = _T_669 | reset; 
  assign _T_672 = _T_671 == 1'h0; 
  assign _T_673 = io_in_a_bits_param == _T_663; 
  assign _T_675 = _T_673 | reset; 
  assign _T_676 = _T_675 == 1'h0; 
  assign _T_677 = io_in_a_bits_size == _T_664; 
  assign _T_679 = _T_677 | reset; 
  assign _T_680 = _T_679 == 1'h0; 
  assign _T_681 = io_in_a_bits_source == _T_665; 
  assign _T_683 = _T_681 | reset; 
  assign _T_684 = _T_683 == 1'h0; 
  assign _T_685 = io_in_a_bits_address == _T_666; 
  assign _T_687 = _T_685 | reset; 
  assign _T_688 = _T_687 == 1'h0; 
  assign _T_690 = _T_642 & _T_654; 
  assign _T_691 = io_in_d_ready & io_in_d_valid; 
  assign _T_693 = 13'h3f << io_in_d_bits_size; 
  assign _T_694 = _T_693[5:0]; 
  assign _T_695 = ~ _T_694; 
  assign _T_696 = _T_695[5:2]; 
  assign _T_697 = io_in_d_bits_opcode[0]; 
  assign _T_701 = _T_699 - 4'h1; 
  assign _T_702 = _T_699 == 4'h0; 
  assign _T_716 = _T_702 == 1'h0; 
  assign _T_717 = io_in_d_valid & _T_716; 
  assign _T_718 = io_in_d_bits_opcode == _T_710; 
  assign _T_720 = _T_718 | reset; 
  assign _T_721 = _T_720 == 1'h0; 
  assign _T_722 = io_in_d_bits_param == _T_711; 
  assign _T_724 = _T_722 | reset; 
  assign _T_725 = _T_724 == 1'h0; 
  assign _T_726 = io_in_d_bits_size == _T_712; 
  assign _T_728 = _T_726 | reset; 
  assign _T_729 = _T_728 == 1'h0; 
  assign _T_730 = io_in_d_bits_source == _T_713; 
  assign _T_732 = _T_730 | reset; 
  assign _T_733 = _T_732 == 1'h0; 
  assign _T_734 = io_in_d_bits_sink == _T_714; 
  assign _T_736 = _T_734 | reset; 
  assign _T_737 = _T_736 == 1'h0; 
  assign _T_738 = io_in_d_bits_denied == _T_715; 
  assign _T_740 = _T_738 | reset; 
  assign _T_741 = _T_740 == 1'h0; 
  assign _T_743 = _T_691 & _T_702; 
  assign _T_756 = _T_754 - 4'h1; 
  assign _T_757 = _T_754 == 4'h0; 
  assign _T_775 = _T_773 - 4'h1; 
  assign _T_776 = _T_773 == 4'h0; 
  assign _T_786 = _T_642 & _T_757; 
  assign _T_788 = 8'h1 << io_in_a_bits_source; 
  assign _T_789 = _T_744 >> io_in_a_bits_source; 
  assign _T_790 = _T_789[0]; 
  assign _T_791 = _T_790 == 1'h0; 
  assign _T_793 = _T_791 | reset; 
  assign _T_794 = _T_793 == 1'h0; 
  assign _GEN_15 = _T_786 ? _T_788 : 8'h0; 
  assign _T_798 = _T_691 & _T_776; 
  assign _T_800 = _T_501 == 1'h0; 
  assign _T_801 = _T_798 & _T_800; 
  assign _T_802 = 8'h1 << io_in_d_bits_source; 
  assign _T_803 = _GEN_15 | _T_744; 
  assign _T_804 = _T_803 >> io_in_d_bits_source; 
  assign _T_805 = _T_804[0]; 
  assign _T_807 = _T_805 | reset; 
  assign _T_808 = _T_807 == 1'h0; 
  assign _GEN_16 = _T_801 ? _T_802 : 8'h0; 
  assign _T_809 = _GEN_15 != _GEN_16; 
  assign _T_810 = _GEN_15 != 8'h0; 
  assign _T_811 = _T_810 == 1'h0; 
  assign _T_812 = _T_809 | _T_811; 
  assign _T_814 = _T_812 | reset; 
  assign _T_815 = _T_814 == 1'h0; 
  assign _T_816 = _T_744 | _GEN_15; 
  assign _T_817 = ~ _GEN_16; 
  assign _T_818 = _T_816 & _T_817; 
  assign _T_820 = _T_744 != 8'h0; 
  assign _T_821 = _T_820 == 1'h0; 
  assign _T_822 = plusarg_reader_out == 32'h0; 
  assign _T_823 = _T_821 | _T_822; 
  assign _T_824 = _T_819 < plusarg_reader_out; 
  assign _T_825 = _T_823 | _T_824; 
  assign _T_827 = _T_825 | reset; 
  assign _T_828 = _T_827 == 1'h0; 
  assign _T_830 = _T_819 + 32'h1; 
  assign _T_833 = _T_642 | _T_691; 
  assign _GEN_19 = io_in_a_valid & _T_96; 
  assign _GEN_35 = io_in_a_valid & _T_154; 
  assign _GEN_53 = io_in_a_valid & _T_216; 
  assign _GEN_65 = io_in_a_valid & _T_261; 
  assign _GEN_75 = io_in_a_valid & _T_302; 
  assign _GEN_85 = io_in_a_valid & _T_345; 
  assign _GEN_95 = io_in_a_valid & _T_391; 
  assign _GEN_105 = io_in_a_valid & _T_437; 
  assign _GEN_115 = io_in_d_valid & _T_501; 
  assign _GEN_125 = io_in_d_valid & _T_521; 
  assign _GEN_137 = io_in_d_valid & _T_549; 
  assign _GEN_149 = io_in_d_valid & _T_578; 
  assign _GEN_155 = io_in_d_valid & _T_595; 
  assign _GEN_161 = io_in_d_valid & _T_613; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_651 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_662 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_663 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_664 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_665 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_666 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_699 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_710 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_711 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_712 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_713 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_714 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_715 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_744 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_754 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_773 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_819 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_651 <= 4'h0;
    end else begin
      if (_T_642) begin
        if (_T_654) begin
          if (_T_649) begin
            _T_651 <= _T_647;
          end else begin
            _T_651 <= 4'h0;
          end
        end else begin
          _T_651 <= _T_653;
        end
      end
    end
    if (_T_690) begin
      _T_662 <= io_in_a_bits_opcode;
    end
    if (_T_690) begin
      _T_663 <= io_in_a_bits_param;
    end
    if (_T_690) begin
      _T_664 <= io_in_a_bits_size;
    end
    if (_T_690) begin
      _T_665 <= io_in_a_bits_source;
    end
    if (_T_690) begin
      _T_666 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_699 <= 4'h0;
    end else begin
      if (_T_691) begin
        if (_T_702) begin
          if (_T_697) begin
            _T_699 <= _T_696;
          end else begin
            _T_699 <= 4'h0;
          end
        end else begin
          _T_699 <= _T_701;
        end
      end
    end
    if (_T_743) begin
      _T_710 <= io_in_d_bits_opcode;
    end
    if (_T_743) begin
      _T_711 <= io_in_d_bits_param;
    end
    if (_T_743) begin
      _T_712 <= io_in_d_bits_size;
    end
    if (_T_743) begin
      _T_713 <= io_in_d_bits_source;
    end
    if (_T_743) begin
      _T_714 <= io_in_d_bits_sink;
    end
    if (_T_743) begin
      _T_715 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_744 <= 8'h0;
    end else begin
      _T_744 <= _T_818;
    end
    if (reset) begin
      _T_754 <= 4'h0;
    end else begin
      if (_T_642) begin
        if (_T_757) begin
          if (_T_649) begin
            _T_754 <= _T_647;
          end else begin
            _T_754 <= 4'h0;
          end
        end else begin
          _T_754 <= _T_756;
        end
      end
    end
    if (reset) begin
      _T_773 <= 4'h0;
    end else begin
      if (_T_691) begin
        if (_T_776) begin
          if (_T_697) begin
            _T_773 <= _T_696;
          end else begin
            _T_773 <= 4'h0;
          end
        end else begin
          _T_773 <= _T_775;
        end
      end
    end
    if (reset) begin
      _T_819 <= 32'h0;
    end else begin
      if (_T_833) begin
        _T_819 <= 32'h0;
      end else begin
        _T_819 <= _T_830;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel has invalid opcode (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:39 assert (TLMessages.isA(bundle.opcode), \"'A' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:46 assert (visible(edge.address(bundle), bundle.source, edge), \"'A' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_127) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_127) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_130) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_130) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_137) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_137) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_140) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_144) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_149) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_149) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_153) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:56 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_153) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_127) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_127) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_130) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_130) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_137) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_137) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_140) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_144) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_206) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_206) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_149) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_149) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_153) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:68 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_153) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_242) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_242) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_140) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_252) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_252) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_256) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_256) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_153) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:77 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_153) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_242) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_242) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_140) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_252) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_252) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_256) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_256) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_242) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_242) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_140) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_252) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_252) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_344) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_344) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_376) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_376) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_140) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_386) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_386) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_256) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_256) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_376) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_376) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_140) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_432) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_432) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_256) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_256) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_242) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_242) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_140) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_140) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_256) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_256) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_153) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:117 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_153) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_481) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_481) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_504) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_504) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_508) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_508) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_512) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_512) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_516) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_516) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_520) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_520) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_504) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_504) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_527) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:285 assert (sink_ok, \"'D' channel Grant carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_527) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_508) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_508) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_535) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_535) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_539) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_539) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_516) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_516) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is denied (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:290 assert (deny_put_ok || !bundle.denied, \"'D' channel Grant is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_504) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_504) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_527) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:295 assert (sink_ok, \"'D' channel GrantData carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_527) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_508) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_508) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_535) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_535) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_539) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_539) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_572) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_572) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:300 assert (deny_get_ok || !bundle.denied, \"'D' channel GrantData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_504) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_504) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_512) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_512) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_516) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_516) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is denied (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:308 assert (deny_put_ok || !bundle.denied, \"'D' channel AccessAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_504) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_504) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_512) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_512) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_572) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_572) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:316 assert (deny_get_ok || !bundle.denied, \"'D' channel AccessAckData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_504) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_504) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_512) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_512) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_516) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_516) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is denied (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:324 assert (deny_put_ok || !bundle.denied, \"'D' channel HintAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel valid and not TL-C (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:341 assert (!bundle.b.valid, \"'B' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel valid and not TL-C (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:342 assert (!bundle.c.valid, \"'C' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel valid and not TL-C (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:343 assert (!bundle.e.valid, \"'E' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_668 & _T_672) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_668 & _T_672) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_668 & _T_676) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_668 & _T_676) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_668 & _T_680) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_668 & _T_680) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_668 & _T_684) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_668 & _T_684) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_668 & _T_688) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_668 & _T_688) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_717 & _T_721) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_717 & _T_721) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_717 & _T_725) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_717 & _T_725) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_717 & _T_729) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_717 & _T_729) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_717 & _T_733) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_717 & _T_733) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_717 & _T_737) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_717 & _T_737) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_717 & _T_741) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_717 & _T_741) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_786 & _T_794) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_786 & _T_794) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_801 & _T_808) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_801 & _T_808) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_815) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_815) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_828) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at ChiplinkTest.scala:220:11)\n    at Monitor.scala:479 assert (!inflight.orR || limit === UInt(0) || watchdog < limit, \"TileLink timeout expired\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_828) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLMonitor_2( 
  input         clock, 
  input         reset, 
  input         io_in_a_ready, 
  input         io_in_a_valid, 
  input  [2:0]  io_in_a_bits_opcode, 
  input  [2:0]  io_in_a_bits_param, 
  input  [2:0]  io_in_a_bits_size, 
  input  [2:0]  io_in_a_bits_source, 
  input  [28:0] io_in_a_bits_address, 
  input  [3:0]  io_in_a_bits_mask, 
  input         io_in_a_bits_corrupt, 
  input         io_in_d_ready, 
  input         io_in_d_valid, 
  input  [2:0]  io_in_d_bits_opcode, 
  input  [1:0]  io_in_d_bits_param, 
  input  [2:0]  io_in_d_bits_size, 
  input  [2:0]  io_in_d_bits_source, 
  input         io_in_d_bits_sink, 
  input         io_in_d_bits_denied, 
  input         io_in_d_bits_corrupt 
);
  wire [31:0] plusarg_reader_out; 
  wire  _T_7; 
  wire  _T_8; 
  wire  _T_22; 
  wire [12:0] _T_24; 
  wire [5:0] _T_25; 
  wire [5:0] _T_26; 
  wire [28:0] _GEN_18; 
  wire [28:0] _T_27; 
  wire  _T_28; 
  wire  _T_30; 
  wire [1:0] _T_31; 
  wire [1:0] _T_33; 
  wire  _T_34; 
  wire  _T_35; 
  wire  _T_36; 
  wire  _T_37; 
  wire  _T_39; 
  wire  _T_40; 
  wire  _T_42; 
  wire  _T_43; 
  wire  _T_44; 
  wire  _T_45; 
  wire  _T_46; 
  wire  _T_47; 
  wire  _T_48; 
  wire  _T_49; 
  wire  _T_50; 
  wire  _T_51; 
  wire  _T_52; 
  wire  _T_53; 
  wire  _T_54; 
  wire  _T_55; 
  wire  _T_56; 
  wire  _T_57; 
  wire  _T_58; 
  wire [3:0] _T_61; 
  wire  _T_96; 
  wire  _T_98; 
  wire [28:0] _T_101; 
  wire [29:0] _T_102; 
  wire [29:0] _T_103; 
  wire [29:0] _T_104; 
  wire  _T_105; 
  wire  _T_106; 
  wire  _T_109; 
  wire  _T_110; 
  wire  _T_113; 
  wire  _T_115; 
  wire  _T_116; 
  wire  _T_119; 
  wire  _T_120; 
  wire  _T_122; 
  wire  _T_123; 
  wire  _T_124; 
  wire  _T_126; 
  wire  _T_127; 
  wire [3:0] _T_128; 
  wire  _T_129; 
  wire  _T_131; 
  wire  _T_132; 
  wire  _T_133; 
  wire  _T_135; 
  wire  _T_136; 
  wire  _T_137; 
  wire  _T_169; 
  wire  _T_171; 
  wire  _T_172; 
  wire  _T_182; 
  wire  _T_203; 
  wire  _T_205; 
  wire  _T_206; 
  wire  _T_207; 
  wire  _T_209; 
  wire  _T_210; 
  wire  _T_215; 
  wire  _T_244; 
  wire [3:0] _T_269; 
  wire [3:0] _T_270; 
  wire  _T_271; 
  wire  _T_273; 
  wire  _T_274; 
  wire  _T_275; 
  wire  _T_296; 
  wire  _T_298; 
  wire  _T_299; 
  wire  _T_304; 
  wire  _T_325; 
  wire  _T_327; 
  wire  _T_328; 
  wire  _T_333; 
  wire  _T_362; 
  wire  _T_364; 
  wire  _T_365; 
  wire  _T_368; 
  wire  _T_369; 
  wire  _T_383; 
  wire  _T_384; 
  wire  _T_385; 
  wire  _T_387; 
  wire  _T_388; 
  wire  _T_389; 
  wire  _T_391; 
  wire  _T_392; 
  wire  _T_393; 
  wire  _T_395; 
  wire  _T_396; 
  wire  _T_397; 
  wire  _T_399; 
  wire  _T_400; 
  wire  _T_401; 
  wire  _T_403; 
  wire  _T_404; 
  wire  _T_405; 
  wire  _T_410; 
  wire  _T_411; 
  wire  _T_416; 
  wire  _T_418; 
  wire  _T_419; 
  wire  _T_420; 
  wire  _T_422; 
  wire  _T_423; 
  wire  _T_433; 
  wire  _T_453; 
  wire  _T_455; 
  wire  _T_456; 
  wire  _T_462; 
  wire  _T_479; 
  wire  _T_497; 
  wire  _T_526; 
  wire [3:0] _T_531; 
  wire  _T_532; 
  wire  _T_533; 
  reg [3:0] _T_535; 
  reg [31:0] _RAND_0;
  wire [3:0] _T_537; 
  wire  _T_538; 
  reg [2:0] _T_546; 
  reg [31:0] _RAND_1;
  reg [2:0] _T_547; 
  reg [31:0] _RAND_2;
  reg [2:0] _T_548; 
  reg [31:0] _RAND_3;
  reg [2:0] _T_549; 
  reg [31:0] _RAND_4;
  reg [28:0] _T_550; 
  reg [31:0] _RAND_5;
  wire  _T_551; 
  wire  _T_552; 
  wire  _T_553; 
  wire  _T_555; 
  wire  _T_556; 
  wire  _T_557; 
  wire  _T_559; 
  wire  _T_560; 
  wire  _T_561; 
  wire  _T_563; 
  wire  _T_564; 
  wire  _T_565; 
  wire  _T_567; 
  wire  _T_568; 
  wire  _T_569; 
  wire  _T_571; 
  wire  _T_572; 
  wire  _T_574; 
  wire  _T_575; 
  wire [12:0] _T_577; 
  wire [5:0] _T_578; 
  wire [5:0] _T_579; 
  wire [3:0] _T_580; 
  wire  _T_581; 
  reg [3:0] _T_583; 
  reg [31:0] _RAND_6;
  wire [3:0] _T_585; 
  wire  _T_586; 
  reg [2:0] _T_594; 
  reg [31:0] _RAND_7;
  reg [1:0] _T_595; 
  reg [31:0] _RAND_8;
  reg [2:0] _T_596; 
  reg [31:0] _RAND_9;
  reg [2:0] _T_597; 
  reg [31:0] _RAND_10;
  reg  _T_598; 
  reg [31:0] _RAND_11;
  reg  _T_599; 
  reg [31:0] _RAND_12;
  wire  _T_600; 
  wire  _T_601; 
  wire  _T_602; 
  wire  _T_604; 
  wire  _T_605; 
  wire  _T_606; 
  wire  _T_608; 
  wire  _T_609; 
  wire  _T_610; 
  wire  _T_612; 
  wire  _T_613; 
  wire  _T_614; 
  wire  _T_616; 
  wire  _T_617; 
  wire  _T_618; 
  wire  _T_620; 
  wire  _T_621; 
  wire  _T_622; 
  wire  _T_624; 
  wire  _T_625; 
  wire  _T_627; 
  reg [7:0] _T_628; 
  reg [31:0] _RAND_13;
  reg [3:0] _T_638; 
  reg [31:0] _RAND_14;
  wire [3:0] _T_640; 
  wire  _T_641; 
  reg [3:0] _T_657; 
  reg [31:0] _RAND_15;
  wire [3:0] _T_659; 
  wire  _T_660; 
  wire  _T_670; 
  wire [7:0] _T_672; 
  wire [7:0] _T_673; 
  wire  _T_674; 
  wire  _T_675; 
  wire  _T_677; 
  wire  _T_678; 
  wire [7:0] _GEN_15; 
  wire  _T_682; 
  wire  _T_684; 
  wire  _T_685; 
  wire [7:0] _T_686; 
  wire [7:0] _T_687; 
  wire [7:0] _T_688; 
  wire  _T_689; 
  wire  _T_691; 
  wire  _T_692; 
  wire [7:0] _GEN_16; 
  wire  _T_693; 
  wire  _T_694; 
  wire  _T_695; 
  wire  _T_696; 
  wire  _T_698; 
  wire  _T_699; 
  wire [7:0] _T_700; 
  wire [7:0] _T_701; 
  wire [7:0] _T_702; 
  reg [31:0] _T_703; 
  reg [31:0] _RAND_16;
  wire  _T_704; 
  wire  _T_705; 
  wire  _T_706; 
  wire  _T_707; 
  wire  _T_708; 
  wire  _T_709; 
  wire  _T_711; 
  wire  _T_712; 
  wire [31:0] _T_714; 
  wire  _T_717; 
  wire  _GEN_19; 
  wire  _GEN_35; 
  wire  _GEN_53; 
  wire  _GEN_65; 
  wire  _GEN_75; 
  wire  _GEN_85; 
  wire  _GEN_95; 
  wire  _GEN_105; 
  wire  _GEN_115; 
  wire  _GEN_125; 
  wire  _GEN_137; 
  wire  _GEN_149; 
  wire  _GEN_155; 
  wire  _GEN_161; 
  dual_plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0)) plusarg_reader ( 
    .out(plusarg_reader_out)
  );
  assign _T_7 = io_in_a_bits_source[2:2]; 
  assign _T_8 = _T_7 == 1'h0; 
  assign _T_22 = _T_8 | _T_7; 
  assign _T_24 = 13'h3f << io_in_a_bits_size; 
  assign _T_25 = _T_24[5:0]; 
  assign _T_26 = ~ _T_25; 
  assign _GEN_18 = {{23'd0}, _T_26}; 
  assign _T_27 = io_in_a_bits_address & _GEN_18; 
  assign _T_28 = _T_27 == 29'h0; 
  assign _T_30 = io_in_a_bits_size[0]; 
  assign _T_31 = 2'h1 << _T_30; 
  assign _T_33 = _T_31 | 2'h1; 
  assign _T_34 = io_in_a_bits_size >= 3'h2; 
  assign _T_35 = _T_33[1]; 
  assign _T_36 = io_in_a_bits_address[1]; 
  assign _T_37 = _T_36 == 1'h0; 
  assign _T_39 = _T_35 & _T_37; 
  assign _T_40 = _T_34 | _T_39; 
  assign _T_42 = _T_35 & _T_36; 
  assign _T_43 = _T_34 | _T_42; 
  assign _T_44 = _T_33[0]; 
  assign _T_45 = io_in_a_bits_address[0]; 
  assign _T_46 = _T_45 == 1'h0; 
  assign _T_47 = _T_37 & _T_46; 
  assign _T_48 = _T_44 & _T_47; 
  assign _T_49 = _T_40 | _T_48; 
  assign _T_50 = _T_37 & _T_45; 
  assign _T_51 = _T_44 & _T_50; 
  assign _T_52 = _T_40 | _T_51; 
  assign _T_53 = _T_36 & _T_46; 
  assign _T_54 = _T_44 & _T_53; 
  assign _T_55 = _T_43 | _T_54; 
  assign _T_56 = _T_36 & _T_45; 
  assign _T_57 = _T_44 & _T_56; 
  assign _T_58 = _T_43 | _T_57; 
  assign _T_61 = {_T_58,_T_55,_T_52,_T_49}; 
  assign _T_96 = io_in_a_bits_opcode == 3'h6; 
  assign _T_98 = io_in_a_bits_size <= 3'h6; 
  assign _T_101 = io_in_a_bits_address ^ 29'h10000000; 
  assign _T_102 = {1'b0,$signed(_T_101)}; 
  assign _T_103 = $signed(_T_102) & $signed(-30'sh10000000); 
  assign _T_104 = $signed(_T_103); 
  assign _T_105 = $signed(_T_104) == $signed(30'sh0); 
  assign _T_106 = _T_98 & _T_105; 
  assign _T_109 = _T_106 | reset; 
  assign _T_110 = _T_109 == 1'h0; 
  assign _T_113 = reset == 1'h0; 
  assign _T_115 = _T_22 | reset; 
  assign _T_116 = _T_115 == 1'h0; 
  assign _T_119 = _T_34 | reset; 
  assign _T_120 = _T_119 == 1'h0; 
  assign _T_122 = _T_28 | reset; 
  assign _T_123 = _T_122 == 1'h0; 
  assign _T_124 = io_in_a_bits_param <= 3'h2; 
  assign _T_126 = _T_124 | reset; 
  assign _T_127 = _T_126 == 1'h0; 
  assign _T_128 = ~ io_in_a_bits_mask; 
  assign _T_129 = _T_128 == 4'h0; 
  assign _T_131 = _T_129 | reset; 
  assign _T_132 = _T_131 == 1'h0; 
  assign _T_133 = io_in_a_bits_corrupt == 1'h0; 
  assign _T_135 = _T_133 | reset; 
  assign _T_136 = _T_135 == 1'h0; 
  assign _T_137 = io_in_a_bits_opcode == 3'h7; 
  assign _T_169 = io_in_a_bits_param != 3'h0; 
  assign _T_171 = _T_169 | reset; 
  assign _T_172 = _T_171 == 1'h0; 
  assign _T_182 = io_in_a_bits_opcode == 3'h4; 
  assign _T_203 = io_in_a_bits_param == 3'h0; 
  assign _T_205 = _T_203 | reset; 
  assign _T_206 = _T_205 == 1'h0; 
  assign _T_207 = io_in_a_bits_mask == _T_61; 
  assign _T_209 = _T_207 | reset; 
  assign _T_210 = _T_209 == 1'h0; 
  assign _T_215 = io_in_a_bits_opcode == 3'h0; 
  assign _T_244 = io_in_a_bits_opcode == 3'h1; 
  assign _T_269 = ~ _T_61; 
  assign _T_270 = io_in_a_bits_mask & _T_269; 
  assign _T_271 = _T_270 == 4'h0; 
  assign _T_273 = _T_271 | reset; 
  assign _T_274 = _T_273 == 1'h0; 
  assign _T_275 = io_in_a_bits_opcode == 3'h2; 
  assign _T_296 = io_in_a_bits_param <= 3'h4; 
  assign _T_298 = _T_296 | reset; 
  assign _T_299 = _T_298 == 1'h0; 
  assign _T_304 = io_in_a_bits_opcode == 3'h3; 
  assign _T_325 = io_in_a_bits_param <= 3'h3; 
  assign _T_327 = _T_325 | reset; 
  assign _T_328 = _T_327 == 1'h0; 
  assign _T_333 = io_in_a_bits_opcode == 3'h5; 
  assign _T_362 = io_in_d_bits_opcode <= 3'h6; 
  assign _T_364 = _T_362 | reset; 
  assign _T_365 = _T_364 == 1'h0; 
  assign _T_368 = io_in_d_bits_source[2:2]; 
  assign _T_369 = _T_368 == 1'h0; 
  assign _T_383 = _T_369 | _T_368; 
  assign _T_384 = io_in_d_bits_sink < 1'h1; 
  assign _T_385 = io_in_d_bits_opcode == 3'h6; 
  assign _T_387 = _T_383 | reset; 
  assign _T_388 = _T_387 == 1'h0; 
  assign _T_389 = io_in_d_bits_size >= 3'h2; 
  assign _T_391 = _T_389 | reset; 
  assign _T_392 = _T_391 == 1'h0; 
  assign _T_393 = io_in_d_bits_param == 2'h0; 
  assign _T_395 = _T_393 | reset; 
  assign _T_396 = _T_395 == 1'h0; 
  assign _T_397 = io_in_d_bits_corrupt == 1'h0; 
  assign _T_399 = _T_397 | reset; 
  assign _T_400 = _T_399 == 1'h0; 
  assign _T_401 = io_in_d_bits_denied == 1'h0; 
  assign _T_403 = _T_401 | reset; 
  assign _T_404 = _T_403 == 1'h0; 
  assign _T_405 = io_in_d_bits_opcode == 3'h4; 
  assign _T_410 = _T_384 | reset; 
  assign _T_411 = _T_410 == 1'h0; 
  assign _T_416 = io_in_d_bits_param <= 2'h2; 
  assign _T_418 = _T_416 | reset; 
  assign _T_419 = _T_418 == 1'h0; 
  assign _T_420 = io_in_d_bits_param != 2'h2; 
  assign _T_422 = _T_420 | reset; 
  assign _T_423 = _T_422 == 1'h0; 
  assign _T_433 = io_in_d_bits_opcode == 3'h5; 
  assign _T_453 = _T_401 | io_in_d_bits_corrupt; 
  assign _T_455 = _T_453 | reset; 
  assign _T_456 = _T_455 == 1'h0; 
  assign _T_462 = io_in_d_bits_opcode == 3'h0; 
  assign _T_479 = io_in_d_bits_opcode == 3'h1; 
  assign _T_497 = io_in_d_bits_opcode == 3'h2; 
  assign _T_526 = io_in_a_ready & io_in_a_valid; 
  assign _T_531 = _T_26[5:2]; 
  assign _T_532 = io_in_a_bits_opcode[2]; 
  assign _T_533 = _T_532 == 1'h0; 
  assign _T_537 = _T_535 - 4'h1; 
  assign _T_538 = _T_535 == 4'h0; 
  assign _T_551 = _T_538 == 1'h0; 
  assign _T_552 = io_in_a_valid & _T_551; 
  assign _T_553 = io_in_a_bits_opcode == _T_546; 
  assign _T_555 = _T_553 | reset; 
  assign _T_556 = _T_555 == 1'h0; 
  assign _T_557 = io_in_a_bits_param == _T_547; 
  assign _T_559 = _T_557 | reset; 
  assign _T_560 = _T_559 == 1'h0; 
  assign _T_561 = io_in_a_bits_size == _T_548; 
  assign _T_563 = _T_561 | reset; 
  assign _T_564 = _T_563 == 1'h0; 
  assign _T_565 = io_in_a_bits_source == _T_549; 
  assign _T_567 = _T_565 | reset; 
  assign _T_568 = _T_567 == 1'h0; 
  assign _T_569 = io_in_a_bits_address == _T_550; 
  assign _T_571 = _T_569 | reset; 
  assign _T_572 = _T_571 == 1'h0; 
  assign _T_574 = _T_526 & _T_538; 
  assign _T_575 = io_in_d_ready & io_in_d_valid; 
  assign _T_577 = 13'h3f << io_in_d_bits_size; 
  assign _T_578 = _T_577[5:0]; 
  assign _T_579 = ~ _T_578; 
  assign _T_580 = _T_579[5:2]; 
  assign _T_581 = io_in_d_bits_opcode[0]; 
  assign _T_585 = _T_583 - 4'h1; 
  assign _T_586 = _T_583 == 4'h0; 
  assign _T_600 = _T_586 == 1'h0; 
  assign _T_601 = io_in_d_valid & _T_600; 
  assign _T_602 = io_in_d_bits_opcode == _T_594; 
  assign _T_604 = _T_602 | reset; 
  assign _T_605 = _T_604 == 1'h0; 
  assign _T_606 = io_in_d_bits_param == _T_595; 
  assign _T_608 = _T_606 | reset; 
  assign _T_609 = _T_608 == 1'h0; 
  assign _T_610 = io_in_d_bits_size == _T_596; 
  assign _T_612 = _T_610 | reset; 
  assign _T_613 = _T_612 == 1'h0; 
  assign _T_614 = io_in_d_bits_source == _T_597; 
  assign _T_616 = _T_614 | reset; 
  assign _T_617 = _T_616 == 1'h0; 
  assign _T_618 = io_in_d_bits_sink == _T_598; 
  assign _T_620 = _T_618 | reset; 
  assign _T_621 = _T_620 == 1'h0; 
  assign _T_622 = io_in_d_bits_denied == _T_599; 
  assign _T_624 = _T_622 | reset; 
  assign _T_625 = _T_624 == 1'h0; 
  assign _T_627 = _T_575 & _T_586; 
  assign _T_640 = _T_638 - 4'h1; 
  assign _T_641 = _T_638 == 4'h0; 
  assign _T_659 = _T_657 - 4'h1; 
  assign _T_660 = _T_657 == 4'h0; 
  assign _T_670 = _T_526 & _T_641; 
  assign _T_672 = 8'h1 << io_in_a_bits_source; 
  assign _T_673 = _T_628 >> io_in_a_bits_source; 
  assign _T_674 = _T_673[0]; 
  assign _T_675 = _T_674 == 1'h0; 
  assign _T_677 = _T_675 | reset; 
  assign _T_678 = _T_677 == 1'h0; 
  assign _GEN_15 = _T_670 ? _T_672 : 8'h0; 
  assign _T_682 = _T_575 & _T_660; 
  assign _T_684 = _T_385 == 1'h0; 
  assign _T_685 = _T_682 & _T_684; 
  assign _T_686 = 8'h1 << io_in_d_bits_source; 
  assign _T_687 = _GEN_15 | _T_628; 
  assign _T_688 = _T_687 >> io_in_d_bits_source; 
  assign _T_689 = _T_688[0]; 
  assign _T_691 = _T_689 | reset; 
  assign _T_692 = _T_691 == 1'h0; 
  assign _GEN_16 = _T_685 ? _T_686 : 8'h0; 
  assign _T_693 = _GEN_15 != _GEN_16; 
  assign _T_694 = _GEN_15 != 8'h0; 
  assign _T_695 = _T_694 == 1'h0; 
  assign _T_696 = _T_693 | _T_695; 
  assign _T_698 = _T_696 | reset; 
  assign _T_699 = _T_698 == 1'h0; 
  assign _T_700 = _T_628 | _GEN_15; 
  assign _T_701 = ~ _GEN_16; 
  assign _T_702 = _T_700 & _T_701; 
  assign _T_704 = _T_628 != 8'h0; 
  assign _T_705 = _T_704 == 1'h0; 
  assign _T_706 = plusarg_reader_out == 32'h0; 
  assign _T_707 = _T_705 | _T_706; 
  assign _T_708 = _T_703 < plusarg_reader_out; 
  assign _T_709 = _T_707 | _T_708; 
  assign _T_711 = _T_709 | reset; 
  assign _T_712 = _T_711 == 1'h0; 
  assign _T_714 = _T_703 + 32'h1; 
  assign _T_717 = _T_526 | _T_575; 
  assign _GEN_19 = io_in_a_valid & _T_96; 
  assign _GEN_35 = io_in_a_valid & _T_137; 
  assign _GEN_53 = io_in_a_valid & _T_182; 
  assign _GEN_65 = io_in_a_valid & _T_215; 
  assign _GEN_75 = io_in_a_valid & _T_244; 
  assign _GEN_85 = io_in_a_valid & _T_275; 
  assign _GEN_95 = io_in_a_valid & _T_304; 
  assign _GEN_105 = io_in_a_valid & _T_333; 
  assign _GEN_115 = io_in_d_valid & _T_385; 
  assign _GEN_125 = io_in_d_valid & _T_405; 
  assign _GEN_137 = io_in_d_valid & _T_433; 
  assign _GEN_149 = io_in_d_valid & _T_462; 
  assign _GEN_155 = io_in_d_valid & _T_479; 
  assign _GEN_161 = io_in_d_valid & _T_497; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_535 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_546 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_547 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_548 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_549 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_550 = _RAND_5[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_583 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_594 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_595 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_596 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_597 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_598 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_599 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_628 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_638 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_657 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_703 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_535 <= 4'h0;
    end else begin
      if (_T_526) begin
        if (_T_538) begin
          if (_T_533) begin
            _T_535 <= _T_531;
          end else begin
            _T_535 <= 4'h0;
          end
        end else begin
          _T_535 <= _T_537;
        end
      end
    end
    if (_T_574) begin
      _T_546 <= io_in_a_bits_opcode;
    end
    if (_T_574) begin
      _T_547 <= io_in_a_bits_param;
    end
    if (_T_574) begin
      _T_548 <= io_in_a_bits_size;
    end
    if (_T_574) begin
      _T_549 <= io_in_a_bits_source;
    end
    if (_T_574) begin
      _T_550 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_583 <= 4'h0;
    end else begin
      if (_T_575) begin
        if (_T_586) begin
          if (_T_581) begin
            _T_583 <= _T_580;
          end else begin
            _T_583 <= 4'h0;
          end
        end else begin
          _T_583 <= _T_585;
        end
      end
    end
    if (_T_627) begin
      _T_594 <= io_in_d_bits_opcode;
    end
    if (_T_627) begin
      _T_595 <= io_in_d_bits_param;
    end
    if (_T_627) begin
      _T_596 <= io_in_d_bits_size;
    end
    if (_T_627) begin
      _T_597 <= io_in_d_bits_source;
    end
    if (_T_627) begin
      _T_598 <= io_in_d_bits_sink;
    end
    if (_T_627) begin
      _T_599 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_628 <= 8'h0;
    end else begin
      _T_628 <= _T_702;
    end
    if (reset) begin
      _T_638 <= 4'h0;
    end else begin
      if (_T_526) begin
        if (_T_641) begin
          if (_T_533) begin
            _T_638 <= _T_531;
          end else begin
            _T_638 <= 4'h0;
          end
        end else begin
          _T_638 <= _T_640;
        end
      end
    end
    if (reset) begin
      _T_657 <= 4'h0;
    end else begin
      if (_T_575) begin
        if (_T_660) begin
          if (_T_581) begin
            _T_657 <= _T_580;
          end else begin
            _T_657 <= 4'h0;
          end
        end else begin
          _T_657 <= _T_659;
        end
      end
    end
    if (reset) begin
      _T_703 <= 32'h0;
    end else begin
      if (_T_717) begin
        _T_703 <= 32'h0;
      end else begin
        _T_703 <= _T_714;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel has invalid opcode (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:39 assert (TLMessages.isA(bundle.opcode), \"'A' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:46 assert (visible(edge.address(bundle), bundle.source, edge), \"'A' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_110) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_113) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_113) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_120) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_120) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_123) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_123) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_127) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_127) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_132) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_132) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_136) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:56 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_136) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_110) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_113) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_113) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_120) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_120) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_123) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_123) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_127) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_127) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_172) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_172) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_132) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_132) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_136) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:68 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_136) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_110) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_123) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_123) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_206) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_206) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_210) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_210) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_136) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:77 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_136) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_110) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_123) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_123) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_206) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_206) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_210) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_210) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_110) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_123) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_123) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_206) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_206) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_274) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_274) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_110) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_123) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_123) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_299) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_299) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_210) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_210) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_110) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_123) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_123) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_328) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_328) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_210) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_210) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_110) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_123) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_123) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_210) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_210) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_136) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:117 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_136) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_365) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_365) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_388) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_388) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_392) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_392) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_396) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_396) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_400) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_400) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_404) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_404) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_388) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_388) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_411) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:285 assert (sink_ok, \"'D' channel Grant carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_411) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_392) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_392) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_419) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_419) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_423) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_423) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_400) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_400) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is denied (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:290 assert (deny_put_ok || !bundle.denied, \"'D' channel Grant is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_388) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_388) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_411) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:295 assert (sink_ok, \"'D' channel GrantData carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_411) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_392) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_392) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_419) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_419) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_423) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_423) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_456) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_456) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:300 assert (deny_get_ok || !bundle.denied, \"'D' channel GrantData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_388) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_388) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_396) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_396) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_400) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_400) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is denied (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:308 assert (deny_put_ok || !bundle.denied, \"'D' channel AccessAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_388) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_388) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_396) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_396) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_456) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_456) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:316 assert (deny_get_ok || !bundle.denied, \"'D' channel AccessAckData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_388) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_388) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_396) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_396) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_400) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_400) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is denied (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:324 assert (deny_put_ok || !bundle.denied, \"'D' channel HintAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel valid and not TL-C (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:341 assert (!bundle.b.valid, \"'B' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel valid and not TL-C (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:342 assert (!bundle.c.valid, \"'C' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel valid and not TL-C (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:343 assert (!bundle.e.valid, \"'E' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_552 & _T_556) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_552 & _T_556) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_552 & _T_560) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_552 & _T_560) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_552 & _T_564) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_552 & _T_564) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_552 & _T_568) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_552 & _T_568) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_552 & _T_572) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_552 & _T_572) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_601 & _T_605) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_601 & _T_605) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_601 & _T_609) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_601 & _T_609) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_601 & _T_613) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_601 & _T_613) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_601 & _T_617) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_601 & _T_617) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_601 & _T_621) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_601 & _T_621) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_601 & _T_625) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_601 & _T_625) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_670 & _T_678) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_670 & _T_678) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_685 & _T_692) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_685 & _T_692) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_699) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_699) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_712) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at ChiplinkTest.scala:143:13)\n    at Monitor.scala:479 assert (!inflight.orR || limit === UInt(0) || watchdog < limit, \"TileLink timeout expired\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_712) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLMonitor_3( 
  input         clock, 
  input         reset, 
  input         io_in_a_ready, 
  input         io_in_a_valid, 
  input  [2:0]  io_in_a_bits_opcode, 
  input  [2:0]  io_in_a_bits_param, 
  input  [2:0]  io_in_a_bits_size, 
  input  [2:0]  io_in_a_bits_source, 
  input  [31:0] io_in_a_bits_address, 
  input  [3:0]  io_in_a_bits_mask, 
  input         io_in_a_bits_corrupt, 
  input         io_in_d_ready, 
  input         io_in_d_valid, 
  input  [2:0]  io_in_d_bits_opcode, 
  input  [1:0]  io_in_d_bits_param, 
  input  [2:0]  io_in_d_bits_size, 
  input  [2:0]  io_in_d_bits_source, 
  input  [4:0]  io_in_d_bits_sink, 
  input         io_in_d_bits_denied, 
  input         io_in_d_bits_corrupt 
);
  wire [31:0] plusarg_reader_out; 
  wire  _T_7; 
  wire  _T_8; 
  wire  _T_22; 
  wire [12:0] _T_24; 
  wire [5:0] _T_25; 
  wire [5:0] _T_26; 
  wire [31:0] _GEN_18; 
  wire [31:0] _T_27; 
  wire  _T_28; 
  wire  _T_30; 
  wire [1:0] _T_31; 
  wire [1:0] _T_33; 
  wire  _T_34; 
  wire  _T_35; 
  wire  _T_36; 
  wire  _T_37; 
  wire  _T_39; 
  wire  _T_40; 
  wire  _T_42; 
  wire  _T_43; 
  wire  _T_44; 
  wire  _T_45; 
  wire  _T_46; 
  wire  _T_47; 
  wire  _T_48; 
  wire  _T_49; 
  wire  _T_50; 
  wire  _T_51; 
  wire  _T_52; 
  wire  _T_53; 
  wire  _T_54; 
  wire  _T_55; 
  wire  _T_56; 
  wire  _T_57; 
  wire  _T_58; 
  wire [3:0] _T_61; 
  wire  _T_96; 
  wire [31:0] _T_98; 
  wire [32:0] _T_99; 
  wire [32:0] _T_100; 
  wire [32:0] _T_101; 
  wire  _T_102; 
  wire  _T_104; 
  wire [31:0] _T_106; 
  wire [32:0] _T_107; 
  wire [32:0] _T_108; 
  wire [32:0] _T_109; 
  wire  _T_110; 
  wire  _T_111; 
  wire  _T_115; 
  wire  _T_116; 
  wire  _T_119; 
  wire  _T_121; 
  wire  _T_122; 
  wire  _T_125; 
  wire  _T_126; 
  wire  _T_128; 
  wire  _T_129; 
  wire  _T_130; 
  wire  _T_132; 
  wire  _T_133; 
  wire [3:0] _T_134; 
  wire  _T_135; 
  wire  _T_137; 
  wire  _T_138; 
  wire  _T_139; 
  wire  _T_141; 
  wire  _T_142; 
  wire  _T_143; 
  wire  _T_181; 
  wire  _T_183; 
  wire  _T_184; 
  wire  _T_194; 
  wire  _T_196; 
  wire  _T_209; 
  wire  _T_210; 
  wire  _T_213; 
  wire  _T_214; 
  wire  _T_221; 
  wire  _T_223; 
  wire  _T_224; 
  wire  _T_225; 
  wire  _T_227; 
  wire  _T_228; 
  wire  _T_233; 
  wire  _T_268; 
  wire [3:0] _T_299; 
  wire [3:0] _T_300; 
  wire  _T_301; 
  wire  _T_303; 
  wire  _T_304; 
  wire  _T_305; 
  wire  _T_307; 
  wire  _T_321; 
  wire  _T_324; 
  wire  _T_325; 
  wire  _T_332; 
  wire  _T_334; 
  wire  _T_335; 
  wire  _T_340; 
  wire  _T_367; 
  wire  _T_369; 
  wire  _T_370; 
  wire  _T_375; 
  wire  _T_410; 
  wire  _T_412; 
  wire  _T_413; 
  wire  _T_416; 
  wire  _T_417; 
  wire  _T_431; 
  wire  _T_432; 
  wire  _T_433; 
  wire  _T_435; 
  wire  _T_436; 
  wire  _T_437; 
  wire  _T_439; 
  wire  _T_440; 
  wire  _T_441; 
  wire  _T_443; 
  wire  _T_444; 
  wire  _T_445; 
  wire  _T_447; 
  wire  _T_448; 
  wire  _T_449; 
  wire  _T_451; 
  wire  _T_452; 
  wire  _T_453; 
  wire  _T_458; 
  wire  _T_459; 
  wire  _T_464; 
  wire  _T_466; 
  wire  _T_467; 
  wire  _T_468; 
  wire  _T_470; 
  wire  _T_471; 
  wire  _T_481; 
  wire  _T_501; 
  wire  _T_503; 
  wire  _T_504; 
  wire  _T_510; 
  wire  _T_527; 
  wire  _T_545; 
  wire  _T_574; 
  wire [3:0] _T_579; 
  wire  _T_580; 
  wire  _T_581; 
  reg [3:0] _T_583; 
  reg [31:0] _RAND_0;
  wire [3:0] _T_585; 
  wire  _T_586; 
  reg [2:0] _T_594; 
  reg [31:0] _RAND_1;
  reg [2:0] _T_595; 
  reg [31:0] _RAND_2;
  reg [2:0] _T_596; 
  reg [31:0] _RAND_3;
  reg [2:0] _T_597; 
  reg [31:0] _RAND_4;
  reg [31:0] _T_598; 
  reg [31:0] _RAND_5;
  wire  _T_599; 
  wire  _T_600; 
  wire  _T_601; 
  wire  _T_603; 
  wire  _T_604; 
  wire  _T_605; 
  wire  _T_607; 
  wire  _T_608; 
  wire  _T_609; 
  wire  _T_611; 
  wire  _T_612; 
  wire  _T_613; 
  wire  _T_615; 
  wire  _T_616; 
  wire  _T_617; 
  wire  _T_619; 
  wire  _T_620; 
  wire  _T_622; 
  wire  _T_623; 
  wire [12:0] _T_625; 
  wire [5:0] _T_626; 
  wire [5:0] _T_627; 
  wire [3:0] _T_628; 
  wire  _T_629; 
  reg [3:0] _T_631; 
  reg [31:0] _RAND_6;
  wire [3:0] _T_633; 
  wire  _T_634; 
  reg [2:0] _T_642; 
  reg [31:0] _RAND_7;
  reg [1:0] _T_643; 
  reg [31:0] _RAND_8;
  reg [2:0] _T_644; 
  reg [31:0] _RAND_9;
  reg [2:0] _T_645; 
  reg [31:0] _RAND_10;
  reg [4:0] _T_646; 
  reg [31:0] _RAND_11;
  reg  _T_647; 
  reg [31:0] _RAND_12;
  wire  _T_648; 
  wire  _T_649; 
  wire  _T_650; 
  wire  _T_652; 
  wire  _T_653; 
  wire  _T_654; 
  wire  _T_656; 
  wire  _T_657; 
  wire  _T_658; 
  wire  _T_660; 
  wire  _T_661; 
  wire  _T_662; 
  wire  _T_664; 
  wire  _T_665; 
  wire  _T_666; 
  wire  _T_668; 
  wire  _T_669; 
  wire  _T_670; 
  wire  _T_672; 
  wire  _T_673; 
  wire  _T_675; 
  reg [7:0] _T_676; 
  reg [31:0] _RAND_13;
  reg [3:0] _T_686; 
  reg [31:0] _RAND_14;
  wire [3:0] _T_688; 
  wire  _T_689; 
  reg [3:0] _T_705; 
  reg [31:0] _RAND_15;
  wire [3:0] _T_707; 
  wire  _T_708; 
  wire  _T_718; 
  wire [7:0] _T_720; 
  wire [7:0] _T_721; 
  wire  _T_722; 
  wire  _T_723; 
  wire  _T_725; 
  wire  _T_726; 
  wire [7:0] _GEN_15; 
  wire  _T_730; 
  wire  _T_732; 
  wire  _T_733; 
  wire [7:0] _T_734; 
  wire [7:0] _T_735; 
  wire [7:0] _T_736; 
  wire  _T_737; 
  wire  _T_739; 
  wire  _T_740; 
  wire [7:0] _GEN_16; 
  wire  _T_741; 
  wire  _T_742; 
  wire  _T_743; 
  wire  _T_744; 
  wire  _T_746; 
  wire  _T_747; 
  wire [7:0] _T_748; 
  wire [7:0] _T_749; 
  wire [7:0] _T_750; 
  reg [31:0] _T_751; 
  reg [31:0] _RAND_16;
  wire  _T_752; 
  wire  _T_753; 
  wire  _T_754; 
  wire  _T_755; 
  wire  _T_756; 
  wire  _T_757; 
  wire  _T_759; 
  wire  _T_760; 
  wire [31:0] _T_762; 
  wire  _T_765; 
  wire  _GEN_19; 
  wire  _GEN_35; 
  wire  _GEN_53; 
  wire  _GEN_65; 
  wire  _GEN_75; 
  wire  _GEN_85; 
  wire  _GEN_95; 
  wire  _GEN_105; 
  wire  _GEN_115; 
  wire  _GEN_125; 
  wire  _GEN_137; 
  wire  _GEN_149; 
  wire  _GEN_155; 
  wire  _GEN_161; 
  dual_plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0)) plusarg_reader ( 
    .out(plusarg_reader_out)
  );
  assign _T_7 = io_in_a_bits_source[2:2]; 
  assign _T_8 = _T_7 == 1'h0; 
  assign _T_22 = _T_8 | _T_7; 
  assign _T_24 = 13'h3f << io_in_a_bits_size; 
  assign _T_25 = _T_24[5:0]; 
  assign _T_26 = ~ _T_25; 
  assign _GEN_18 = {{26'd0}, _T_26}; 
  assign _T_27 = io_in_a_bits_address & _GEN_18; 
  assign _T_28 = _T_27 == 32'h0; 
  assign _T_30 = io_in_a_bits_size[0]; 
  assign _T_31 = 2'h1 << _T_30; 
  assign _T_33 = _T_31 | 2'h1; 
  assign _T_34 = io_in_a_bits_size >= 3'h2; 
  assign _T_35 = _T_33[1]; 
  assign _T_36 = io_in_a_bits_address[1]; 
  assign _T_37 = _T_36 == 1'h0; 
  assign _T_39 = _T_35 & _T_37; 
  assign _T_40 = _T_34 | _T_39; 
  assign _T_42 = _T_35 & _T_36; 
  assign _T_43 = _T_34 | _T_42; 
  assign _T_44 = _T_33[0]; 
  assign _T_45 = io_in_a_bits_address[0]; 
  assign _T_46 = _T_45 == 1'h0; 
  assign _T_47 = _T_37 & _T_46; 
  assign _T_48 = _T_44 & _T_47; 
  assign _T_49 = _T_40 | _T_48; 
  assign _T_50 = _T_37 & _T_45; 
  assign _T_51 = _T_44 & _T_50; 
  assign _T_52 = _T_40 | _T_51; 
  assign _T_53 = _T_36 & _T_46; 
  assign _T_54 = _T_44 & _T_53; 
  assign _T_55 = _T_43 | _T_54; 
  assign _T_56 = _T_36 & _T_45; 
  assign _T_57 = _T_44 & _T_56; 
  assign _T_58 = _T_43 | _T_57; 
  assign _T_61 = {_T_58,_T_55,_T_52,_T_49}; 
  assign _T_96 = io_in_a_bits_opcode == 3'h6; 
  assign _T_98 = io_in_a_bits_address ^ 32'h40000000; 
  assign _T_99 = {1'b0,$signed(_T_98)}; 
  assign _T_100 = $signed(_T_99) & $signed(-33'sh20000000); 
  assign _T_101 = $signed(_T_100); 
  assign _T_102 = $signed(_T_101) == $signed(33'sh0); 
  assign _T_104 = 3'h6 == io_in_a_bits_size; 
  assign _T_106 = io_in_a_bits_address ^ 32'h80000000; 
  assign _T_107 = {1'b0,$signed(_T_106)}; 
  assign _T_108 = $signed(_T_107) & $signed(-33'sh80000000); 
  assign _T_109 = $signed(_T_108); 
  assign _T_110 = $signed(_T_109) == $signed(33'sh0); 
  assign _T_111 = _T_104 & _T_110; 
  assign _T_115 = _T_111 | reset; 
  assign _T_116 = _T_115 == 1'h0; 
  assign _T_119 = reset == 1'h0; 
  assign _T_121 = _T_22 | reset; 
  assign _T_122 = _T_121 == 1'h0; 
  assign _T_125 = _T_34 | reset; 
  assign _T_126 = _T_125 == 1'h0; 
  assign _T_128 = _T_28 | reset; 
  assign _T_129 = _T_128 == 1'h0; 
  assign _T_130 = io_in_a_bits_param <= 3'h2; 
  assign _T_132 = _T_130 | reset; 
  assign _T_133 = _T_132 == 1'h0; 
  assign _T_134 = ~ io_in_a_bits_mask; 
  assign _T_135 = _T_134 == 4'h0; 
  assign _T_137 = _T_135 | reset; 
  assign _T_138 = _T_137 == 1'h0; 
  assign _T_139 = io_in_a_bits_corrupt == 1'h0; 
  assign _T_141 = _T_139 | reset; 
  assign _T_142 = _T_141 == 1'h0; 
  assign _T_143 = io_in_a_bits_opcode == 3'h7; 
  assign _T_181 = io_in_a_bits_param != 3'h0; 
  assign _T_183 = _T_181 | reset; 
  assign _T_184 = _T_183 == 1'h0; 
  assign _T_194 = io_in_a_bits_opcode == 3'h4; 
  assign _T_196 = io_in_a_bits_size <= 3'h6; 
  assign _T_209 = _T_102 | _T_110; 
  assign _T_210 = _T_196 & _T_209; 
  assign _T_213 = _T_210 | reset; 
  assign _T_214 = _T_213 == 1'h0; 
  assign _T_221 = io_in_a_bits_param == 3'h0; 
  assign _T_223 = _T_221 | reset; 
  assign _T_224 = _T_223 == 1'h0; 
  assign _T_225 = io_in_a_bits_mask == _T_61; 
  assign _T_227 = _T_225 | reset; 
  assign _T_228 = _T_227 == 1'h0; 
  assign _T_233 = io_in_a_bits_opcode == 3'h0; 
  assign _T_268 = io_in_a_bits_opcode == 3'h1; 
  assign _T_299 = ~ _T_61; 
  assign _T_300 = io_in_a_bits_mask & _T_299; 
  assign _T_301 = _T_300 == 4'h0; 
  assign _T_303 = _T_301 | reset; 
  assign _T_304 = _T_303 == 1'h0; 
  assign _T_305 = io_in_a_bits_opcode == 3'h2; 
  assign _T_307 = io_in_a_bits_size <= 3'h3; 
  assign _T_321 = _T_307 & _T_209; 
  assign _T_324 = _T_321 | reset; 
  assign _T_325 = _T_324 == 1'h0; 
  assign _T_332 = io_in_a_bits_param <= 3'h4; 
  assign _T_334 = _T_332 | reset; 
  assign _T_335 = _T_334 == 1'h0; 
  assign _T_340 = io_in_a_bits_opcode == 3'h3; 
  assign _T_367 = io_in_a_bits_param <= 3'h3; 
  assign _T_369 = _T_367 | reset; 
  assign _T_370 = _T_369 == 1'h0; 
  assign _T_375 = io_in_a_bits_opcode == 3'h5; 
  assign _T_410 = io_in_d_bits_opcode <= 3'h6; 
  assign _T_412 = _T_410 | reset; 
  assign _T_413 = _T_412 == 1'h0; 
  assign _T_416 = io_in_d_bits_source[2:2]; 
  assign _T_417 = _T_416 == 1'h0; 
  assign _T_431 = _T_417 | _T_416; 
  assign _T_432 = io_in_d_bits_sink < 5'h1f; 
  assign _T_433 = io_in_d_bits_opcode == 3'h6; 
  assign _T_435 = _T_431 | reset; 
  assign _T_436 = _T_435 == 1'h0; 
  assign _T_437 = io_in_d_bits_size >= 3'h2; 
  assign _T_439 = _T_437 | reset; 
  assign _T_440 = _T_439 == 1'h0; 
  assign _T_441 = io_in_d_bits_param == 2'h0; 
  assign _T_443 = _T_441 | reset; 
  assign _T_444 = _T_443 == 1'h0; 
  assign _T_445 = io_in_d_bits_corrupt == 1'h0; 
  assign _T_447 = _T_445 | reset; 
  assign _T_448 = _T_447 == 1'h0; 
  assign _T_449 = io_in_d_bits_denied == 1'h0; 
  assign _T_451 = _T_449 | reset; 
  assign _T_452 = _T_451 == 1'h0; 
  assign _T_453 = io_in_d_bits_opcode == 3'h4; 
  assign _T_458 = _T_432 | reset; 
  assign _T_459 = _T_458 == 1'h0; 
  assign _T_464 = io_in_d_bits_param <= 2'h2; 
  assign _T_466 = _T_464 | reset; 
  assign _T_467 = _T_466 == 1'h0; 
  assign _T_468 = io_in_d_bits_param != 2'h2; 
  assign _T_470 = _T_468 | reset; 
  assign _T_471 = _T_470 == 1'h0; 
  assign _T_481 = io_in_d_bits_opcode == 3'h5; 
  assign _T_501 = _T_449 | io_in_d_bits_corrupt; 
  assign _T_503 = _T_501 | reset; 
  assign _T_504 = _T_503 == 1'h0; 
  assign _T_510 = io_in_d_bits_opcode == 3'h0; 
  assign _T_527 = io_in_d_bits_opcode == 3'h1; 
  assign _T_545 = io_in_d_bits_opcode == 3'h2; 
  assign _T_574 = io_in_a_ready & io_in_a_valid; 
  assign _T_579 = _T_26[5:2]; 
  assign _T_580 = io_in_a_bits_opcode[2]; 
  assign _T_581 = _T_580 == 1'h0; 
  assign _T_585 = _T_583 - 4'h1; 
  assign _T_586 = _T_583 == 4'h0; 
  assign _T_599 = _T_586 == 1'h0; 
  assign _T_600 = io_in_a_valid & _T_599; 
  assign _T_601 = io_in_a_bits_opcode == _T_594; 
  assign _T_603 = _T_601 | reset; 
  assign _T_604 = _T_603 == 1'h0; 
  assign _T_605 = io_in_a_bits_param == _T_595; 
  assign _T_607 = _T_605 | reset; 
  assign _T_608 = _T_607 == 1'h0; 
  assign _T_609 = io_in_a_bits_size == _T_596; 
  assign _T_611 = _T_609 | reset; 
  assign _T_612 = _T_611 == 1'h0; 
  assign _T_613 = io_in_a_bits_source == _T_597; 
  assign _T_615 = _T_613 | reset; 
  assign _T_616 = _T_615 == 1'h0; 
  assign _T_617 = io_in_a_bits_address == _T_598; 
  assign _T_619 = _T_617 | reset; 
  assign _T_620 = _T_619 == 1'h0; 
  assign _T_622 = _T_574 & _T_586; 
  assign _T_623 = io_in_d_ready & io_in_d_valid; 
  assign _T_625 = 13'h3f << io_in_d_bits_size; 
  assign _T_626 = _T_625[5:0]; 
  assign _T_627 = ~ _T_626; 
  assign _T_628 = _T_627[5:2]; 
  assign _T_629 = io_in_d_bits_opcode[0]; 
  assign _T_633 = _T_631 - 4'h1; 
  assign _T_634 = _T_631 == 4'h0; 
  assign _T_648 = _T_634 == 1'h0; 
  assign _T_649 = io_in_d_valid & _T_648; 
  assign _T_650 = io_in_d_bits_opcode == _T_642; 
  assign _T_652 = _T_650 | reset; 
  assign _T_653 = _T_652 == 1'h0; 
  assign _T_654 = io_in_d_bits_param == _T_643; 
  assign _T_656 = _T_654 | reset; 
  assign _T_657 = _T_656 == 1'h0; 
  assign _T_658 = io_in_d_bits_size == _T_644; 
  assign _T_660 = _T_658 | reset; 
  assign _T_661 = _T_660 == 1'h0; 
  assign _T_662 = io_in_d_bits_source == _T_645; 
  assign _T_664 = _T_662 | reset; 
  assign _T_665 = _T_664 == 1'h0; 
  assign _T_666 = io_in_d_bits_sink == _T_646; 
  assign _T_668 = _T_666 | reset; 
  assign _T_669 = _T_668 == 1'h0; 
  assign _T_670 = io_in_d_bits_denied == _T_647; 
  assign _T_672 = _T_670 | reset; 
  assign _T_673 = _T_672 == 1'h0; 
  assign _T_675 = _T_623 & _T_634; 
  assign _T_688 = _T_686 - 4'h1; 
  assign _T_689 = _T_686 == 4'h0; 
  assign _T_707 = _T_705 - 4'h1; 
  assign _T_708 = _T_705 == 4'h0; 
  assign _T_718 = _T_574 & _T_689; 
  assign _T_720 = 8'h1 << io_in_a_bits_source; 
  assign _T_721 = _T_676 >> io_in_a_bits_source; 
  assign _T_722 = _T_721[0]; 
  assign _T_723 = _T_722 == 1'h0; 
  assign _T_725 = _T_723 | reset; 
  assign _T_726 = _T_725 == 1'h0; 
  assign _GEN_15 = _T_718 ? _T_720 : 8'h0; 
  assign _T_730 = _T_623 & _T_708; 
  assign _T_732 = _T_433 == 1'h0; 
  assign _T_733 = _T_730 & _T_732; 
  assign _T_734 = 8'h1 << io_in_d_bits_source; 
  assign _T_735 = _GEN_15 | _T_676; 
  assign _T_736 = _T_735 >> io_in_d_bits_source; 
  assign _T_737 = _T_736[0]; 
  assign _T_739 = _T_737 | reset; 
  assign _T_740 = _T_739 == 1'h0; 
  assign _GEN_16 = _T_733 ? _T_734 : 8'h0; 
  assign _T_741 = _GEN_15 != _GEN_16; 
  assign _T_742 = _GEN_15 != 8'h0; 
  assign _T_743 = _T_742 == 1'h0; 
  assign _T_744 = _T_741 | _T_743; 
  assign _T_746 = _T_744 | reset; 
  assign _T_747 = _T_746 == 1'h0; 
  assign _T_748 = _T_676 | _GEN_15; 
  assign _T_749 = ~ _GEN_16; 
  assign _T_750 = _T_748 & _T_749; 
  assign _T_752 = _T_676 != 8'h0; 
  assign _T_753 = _T_752 == 1'h0; 
  assign _T_754 = plusarg_reader_out == 32'h0; 
  assign _T_755 = _T_753 | _T_754; 
  assign _T_756 = _T_751 < plusarg_reader_out; 
  assign _T_757 = _T_755 | _T_756; 
  assign _T_759 = _T_757 | reset; 
  assign _T_760 = _T_759 == 1'h0; 
  assign _T_762 = _T_751 + 32'h1; 
  assign _T_765 = _T_574 | _T_623; 
  assign _GEN_19 = io_in_a_valid & _T_96; 
  assign _GEN_35 = io_in_a_valid & _T_143; 
  assign _GEN_53 = io_in_a_valid & _T_194; 
  assign _GEN_65 = io_in_a_valid & _T_233; 
  assign _GEN_75 = io_in_a_valid & _T_268; 
  assign _GEN_85 = io_in_a_valid & _T_305; 
  assign _GEN_95 = io_in_a_valid & _T_340; 
  assign _GEN_105 = io_in_a_valid & _T_375; 
  assign _GEN_115 = io_in_d_valid & _T_433; 
  assign _GEN_125 = io_in_d_valid & _T_453; 
  assign _GEN_137 = io_in_d_valid & _T_481; 
  assign _GEN_149 = io_in_d_valid & _T_510; 
  assign _GEN_155 = io_in_d_valid & _T_527; 
  assign _GEN_161 = io_in_d_valid & _T_545; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_583 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_594 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_595 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_596 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_597 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_598 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_631 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_642 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_643 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_644 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_645 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_646 = _RAND_11[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_647 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_676 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_686 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_705 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_751 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_583 <= 4'h0;
    end else begin
      if (_T_574) begin
        if (_T_586) begin
          if (_T_581) begin
            _T_583 <= _T_579;
          end else begin
            _T_583 <= 4'h0;
          end
        end else begin
          _T_583 <= _T_585;
        end
      end
    end
    if (_T_622) begin
      _T_594 <= io_in_a_bits_opcode;
    end
    if (_T_622) begin
      _T_595 <= io_in_a_bits_param;
    end
    if (_T_622) begin
      _T_596 <= io_in_a_bits_size;
    end
    if (_T_622) begin
      _T_597 <= io_in_a_bits_source;
    end
    if (_T_622) begin
      _T_598 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_631 <= 4'h0;
    end else begin
      if (_T_623) begin
        if (_T_634) begin
          if (_T_629) begin
            _T_631 <= _T_628;
          end else begin
            _T_631 <= 4'h0;
          end
        end else begin
          _T_631 <= _T_633;
        end
      end
    end
    if (_T_675) begin
      _T_642 <= io_in_d_bits_opcode;
    end
    if (_T_675) begin
      _T_643 <= io_in_d_bits_param;
    end
    if (_T_675) begin
      _T_644 <= io_in_d_bits_size;
    end
    if (_T_675) begin
      _T_645 <= io_in_d_bits_source;
    end
    if (_T_675) begin
      _T_646 <= io_in_d_bits_sink;
    end
    if (_T_675) begin
      _T_647 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_676 <= 8'h0;
    end else begin
      _T_676 <= _T_750;
    end
    if (reset) begin
      _T_686 <= 4'h0;
    end else begin
      if (_T_574) begin
        if (_T_689) begin
          if (_T_581) begin
            _T_686 <= _T_579;
          end else begin
            _T_686 <= 4'h0;
          end
        end else begin
          _T_686 <= _T_688;
        end
      end
    end
    if (reset) begin
      _T_705 <= 4'h0;
    end else begin
      if (_T_623) begin
        if (_T_708) begin
          if (_T_629) begin
            _T_705 <= _T_628;
          end else begin
            _T_705 <= 4'h0;
          end
        end else begin
          _T_705 <= _T_707;
        end
      end
    end
    if (reset) begin
      _T_751 <= 32'h0;
    end else begin
      if (_T_765) begin
        _T_751 <= 32'h0;
      end else begin
        _T_751 <= _T_762;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel has invalid opcode (connected at BusBypass.scala:31:12)\n    at Monitor.scala:39 assert (TLMessages.isA(bundle.opcode), \"'A' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:46 assert (visible(edge.address(bundle), bundle.source, edge), \"'A' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at BusBypass.scala:31:12)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_119) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at BusBypass.scala:31:12)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_119) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_122) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at BusBypass.scala:31:12)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_122) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_126) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at BusBypass.scala:31:12)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_126) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at BusBypass.scala:31:12)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_129) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at BusBypass.scala:31:12)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_138) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at BusBypass.scala:31:12)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_138) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_142) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at BusBypass.scala:31:12)\n    at Monitor.scala:56 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_142) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at BusBypass.scala:31:12)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_119) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at BusBypass.scala:31:12)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_119) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_122) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at BusBypass.scala:31:12)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_122) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_126) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at BusBypass.scala:31:12)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_126) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at BusBypass.scala:31:12)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_129) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at BusBypass.scala:31:12)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_184) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at BusBypass.scala:31:12)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_184) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_138) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at BusBypass.scala:31:12)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_138) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_142) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at BusBypass.scala:31:12)\n    at Monitor.scala:68 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_142) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_214) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at BusBypass.scala:31:12)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_214) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_122) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at BusBypass.scala:31:12)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_122) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at BusBypass.scala:31:12)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_129) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_224) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at BusBypass.scala:31:12)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_224) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_228) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at BusBypass.scala:31:12)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_228) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_142) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at BusBypass.scala:31:12)\n    at Monitor.scala:77 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_142) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_214) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at BusBypass.scala:31:12)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_214) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_122) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at BusBypass.scala:31:12)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_122) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at BusBypass.scala:31:12)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_129) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_224) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at BusBypass.scala:31:12)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_224) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_228) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at BusBypass.scala:31:12)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_228) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_214) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at BusBypass.scala:31:12)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_214) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_122) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at BusBypass.scala:31:12)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_122) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at BusBypass.scala:31:12)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_129) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_224) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at BusBypass.scala:31:12)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_224) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_304) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at BusBypass.scala:31:12)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_304) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_325) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at BusBypass.scala:31:12)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_325) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_122) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at BusBypass.scala:31:12)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_122) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at BusBypass.scala:31:12)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_129) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_335) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at BusBypass.scala:31:12)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_335) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_228) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at BusBypass.scala:31:12)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_228) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_325) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at BusBypass.scala:31:12)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_325) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_122) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at BusBypass.scala:31:12)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_122) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at BusBypass.scala:31:12)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_129) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_370) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at BusBypass.scala:31:12)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_370) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_228) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at BusBypass.scala:31:12)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_228) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_214) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at BusBypass.scala:31:12)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_214) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_122) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at BusBypass.scala:31:12)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_122) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at BusBypass.scala:31:12)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_129) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_228) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at BusBypass.scala:31:12)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_228) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_142) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at BusBypass.scala:31:12)\n    at Monitor.scala:117 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_142) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_413) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at BusBypass.scala:31:12)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_413) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_436) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at BusBypass.scala:31:12)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_436) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_440) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at BusBypass.scala:31:12)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_440) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_444) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at BusBypass.scala:31:12)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_444) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_448) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at BusBypass.scala:31:12)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_448) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_452) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at BusBypass.scala:31:12)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_452) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_436) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at BusBypass.scala:31:12)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_436) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_459) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at BusBypass.scala:31:12)\n    at Monitor.scala:285 assert (sink_ok, \"'D' channel Grant carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_459) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_440) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at BusBypass.scala:31:12)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_440) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_467) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at BusBypass.scala:31:12)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_467) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_471) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at BusBypass.scala:31:12)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_471) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_448) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at BusBypass.scala:31:12)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_448) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is denied (connected at BusBypass.scala:31:12)\n    at Monitor.scala:290 assert (deny_put_ok || !bundle.denied, \"'D' channel Grant is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_436) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at BusBypass.scala:31:12)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_436) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_459) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at BusBypass.scala:31:12)\n    at Monitor.scala:295 assert (sink_ok, \"'D' channel GrantData carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_459) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_440) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at BusBypass.scala:31:12)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_440) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_467) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at BusBypass.scala:31:12)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_467) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_471) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at BusBypass.scala:31:12)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_471) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_504) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at BusBypass.scala:31:12)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_504) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied (connected at BusBypass.scala:31:12)\n    at Monitor.scala:300 assert (deny_get_ok || !bundle.denied, \"'D' channel GrantData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_436) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at BusBypass.scala:31:12)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_436) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_444) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at BusBypass.scala:31:12)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_444) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_448) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at BusBypass.scala:31:12)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_448) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is denied (connected at BusBypass.scala:31:12)\n    at Monitor.scala:308 assert (deny_put_ok || !bundle.denied, \"'D' channel AccessAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_436) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at BusBypass.scala:31:12)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_436) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_444) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at BusBypass.scala:31:12)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_444) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_504) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at BusBypass.scala:31:12)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_504) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied (connected at BusBypass.scala:31:12)\n    at Monitor.scala:316 assert (deny_get_ok || !bundle.denied, \"'D' channel AccessAckData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_436) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at BusBypass.scala:31:12)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_436) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_444) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at BusBypass.scala:31:12)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_444) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_448) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at BusBypass.scala:31:12)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_448) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is denied (connected at BusBypass.scala:31:12)\n    at Monitor.scala:324 assert (deny_put_ok || !bundle.denied, \"'D' channel HintAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel valid and not TL-C (connected at BusBypass.scala:31:12)\n    at Monitor.scala:341 assert (!bundle.b.valid, \"'B' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel valid and not TL-C (connected at BusBypass.scala:31:12)\n    at Monitor.scala:342 assert (!bundle.c.valid, \"'C' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel valid and not TL-C (connected at BusBypass.scala:31:12)\n    at Monitor.scala:343 assert (!bundle.e.valid, \"'E' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_600 & _T_604) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at BusBypass.scala:31:12)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_600 & _T_604) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_600 & _T_608) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at BusBypass.scala:31:12)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_600 & _T_608) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_600 & _T_612) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at BusBypass.scala:31:12)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_600 & _T_612) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_600 & _T_616) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at BusBypass.scala:31:12)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_600 & _T_616) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_600 & _T_620) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at BusBypass.scala:31:12)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_600 & _T_620) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_649 & _T_653) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at BusBypass.scala:31:12)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_649 & _T_653) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_649 & _T_657) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at BusBypass.scala:31:12)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_649 & _T_657) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_649 & _T_661) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at BusBypass.scala:31:12)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_649 & _T_661) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_649 & _T_665) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at BusBypass.scala:31:12)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_649 & _T_665) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_649 & _T_669) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at BusBypass.scala:31:12)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_649 & _T_669) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_649 & _T_673) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at BusBypass.scala:31:12)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_649 & _T_673) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_718 & _T_726) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at BusBypass.scala:31:12)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_718 & _T_726) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_733 & _T_740) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at BusBypass.scala:31:12)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_733 & _T_740) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_747) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 8 (connected at BusBypass.scala:31:12)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_747) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_760) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at BusBypass.scala:31:12)\n    at Monitor.scala:479 assert (!inflight.orR || limit === UInt(0) || watchdog < limit, \"TileLink timeout expired\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_760) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLMonitor_4( 
  input          clock, 
  input          reset, 
  input          io_in_a_ready, 
  input          io_in_a_valid, 
  input  [2:0]   io_in_a_bits_opcode, 
  input  [2:0]   io_in_a_bits_param, 
  input  [3:0]   io_in_a_bits_size, 
  input  [2:0]   io_in_a_bits_source, 
  input  [127:0] io_in_a_bits_address, 
  input  [3:0]   io_in_a_bits_mask, 
  input          io_in_a_bits_corrupt, 
  input          io_in_d_ready, 
  input          io_in_d_valid, 
  input  [2:0]   io_in_d_bits_opcode, 
  input  [1:0]   io_in_d_bits_param, 
  input  [3:0]   io_in_d_bits_size, 
  input  [2:0]   io_in_d_bits_source, 
  input          io_in_d_bits_sink, 
  input          io_in_d_bits_denied, 
  input          io_in_d_bits_corrupt 
);
  wire [31:0] plusarg_reader_out; 
  wire  _T_7; 
  wire  _T_8; 
  wire  _T_22; 
  wire [26:0] _T_24; 
  wire [11:0] _T_25; 
  wire [11:0] _T_26; 
  wire [127:0] _GEN_18; 
  wire [127:0] _T_27; 
  wire  _T_28; 
  wire  _T_30; 
  wire [1:0] _T_31; 
  wire [1:0] _T_33; 
  wire  _T_34; 
  wire  _T_35; 
  wire  _T_36; 
  wire  _T_37; 
  wire  _T_39; 
  wire  _T_40; 
  wire  _T_42; 
  wire  _T_43; 
  wire  _T_44; 
  wire  _T_45; 
  wire  _T_46; 
  wire  _T_47; 
  wire  _T_48; 
  wire  _T_49; 
  wire  _T_50; 
  wire  _T_51; 
  wire  _T_52; 
  wire  _T_53; 
  wire  _T_54; 
  wire  _T_55; 
  wire  _T_56; 
  wire  _T_57; 
  wire  _T_58; 
  wire [3:0] _T_61; 
  wire [128:0] _T_72; 
  wire  _T_96; 
  wire  _T_98; 
  wire [128:0] _T_103; 
  wire [128:0] _T_104; 
  wire  _T_105; 
  wire  _T_106; 
  wire  _T_109; 
  wire  _T_110; 
  wire  _T_113; 
  wire  _T_115; 
  wire  _T_116; 
  wire  _T_119; 
  wire  _T_120; 
  wire  _T_122; 
  wire  _T_123; 
  wire  _T_124; 
  wire  _T_126; 
  wire  _T_127; 
  wire [3:0] _T_128; 
  wire  _T_129; 
  wire  _T_131; 
  wire  _T_132; 
  wire  _T_133; 
  wire  _T_135; 
  wire  _T_136; 
  wire  _T_137; 
  wire  _T_169; 
  wire  _T_171; 
  wire  _T_172; 
  wire  _T_182; 
  wire  _T_203; 
  wire  _T_205; 
  wire  _T_206; 
  wire  _T_207; 
  wire  _T_209; 
  wire  _T_210; 
  wire  _T_215; 
  wire  _T_244; 
  wire [3:0] _T_269; 
  wire [3:0] _T_270; 
  wire  _T_271; 
  wire  _T_273; 
  wire  _T_274; 
  wire  _T_275; 
  wire  _T_277; 
  wire  _T_285; 
  wire  _T_288; 
  wire  _T_289; 
  wire  _T_296; 
  wire  _T_298; 
  wire  _T_299; 
  wire  _T_304; 
  wire  _T_325; 
  wire  _T_327; 
  wire  _T_328; 
  wire  _T_333; 
  wire  _T_362; 
  wire  _T_364; 
  wire  _T_365; 
  wire  _T_368; 
  wire  _T_369; 
  wire  _T_383; 
  wire  _T_384; 
  wire  _T_385; 
  wire  _T_387; 
  wire  _T_388; 
  wire  _T_389; 
  wire  _T_391; 
  wire  _T_392; 
  wire  _T_393; 
  wire  _T_395; 
  wire  _T_396; 
  wire  _T_397; 
  wire  _T_399; 
  wire  _T_400; 
  wire  _T_401; 
  wire  _T_403; 
  wire  _T_404; 
  wire  _T_405; 
  wire  _T_410; 
  wire  _T_411; 
  wire  _T_416; 
  wire  _T_418; 
  wire  _T_419; 
  wire  _T_420; 
  wire  _T_422; 
  wire  _T_423; 
  wire  _T_433; 
  wire  _T_453; 
  wire  _T_455; 
  wire  _T_456; 
  wire  _T_462; 
  wire  _T_479; 
  wire  _T_497; 
  wire  _T_526; 
  wire [9:0] _T_531; 
  wire  _T_532; 
  wire  _T_533; 
  reg [9:0] _T_535; 
  reg [31:0] _RAND_0;
  wire [9:0] _T_537; 
  wire  _T_538; 
  reg [2:0] _T_546; 
  reg [31:0] _RAND_1;
  reg [2:0] _T_547; 
  reg [31:0] _RAND_2;
  reg [3:0] _T_548; 
  reg [31:0] _RAND_3;
  reg [2:0] _T_549; 
  reg [31:0] _RAND_4;
  reg [127:0] _T_550; 
  reg [127:0] _RAND_5;
  wire  _T_551; 
  wire  _T_552; 
  wire  _T_553; 
  wire  _T_555; 
  wire  _T_556; 
  wire  _T_557; 
  wire  _T_559; 
  wire  _T_560; 
  wire  _T_561; 
  wire  _T_563; 
  wire  _T_564; 
  wire  _T_565; 
  wire  _T_567; 
  wire  _T_568; 
  wire  _T_569; 
  wire  _T_571; 
  wire  _T_572; 
  wire  _T_574; 
  wire  _T_575; 
  wire [26:0] _T_577; 
  wire [11:0] _T_578; 
  wire [11:0] _T_579; 
  wire [9:0] _T_580; 
  wire  _T_581; 
  reg [9:0] _T_583; 
  reg [31:0] _RAND_6;
  wire [9:0] _T_585; 
  wire  _T_586; 
  reg [2:0] _T_594; 
  reg [31:0] _RAND_7;
  reg [1:0] _T_595; 
  reg [31:0] _RAND_8;
  reg [3:0] _T_596; 
  reg [31:0] _RAND_9;
  reg [2:0] _T_597; 
  reg [31:0] _RAND_10;
  reg  _T_598; 
  reg [31:0] _RAND_11;
  reg  _T_599; 
  reg [31:0] _RAND_12;
  wire  _T_600; 
  wire  _T_601; 
  wire  _T_602; 
  wire  _T_604; 
  wire  _T_605; 
  wire  _T_606; 
  wire  _T_608; 
  wire  _T_609; 
  wire  _T_610; 
  wire  _T_612; 
  wire  _T_613; 
  wire  _T_614; 
  wire  _T_616; 
  wire  _T_617; 
  wire  _T_618; 
  wire  _T_620; 
  wire  _T_621; 
  wire  _T_622; 
  wire  _T_624; 
  wire  _T_625; 
  wire  _T_627; 
  reg [7:0] _T_628; 
  reg [31:0] _RAND_13;
  reg [9:0] _T_638; 
  reg [31:0] _RAND_14;
  wire [9:0] _T_640; 
  wire  _T_641; 
  reg [9:0] _T_657; 
  reg [31:0] _RAND_15;
  wire [9:0] _T_659; 
  wire  _T_660; 
  wire  _T_670; 
  wire [7:0] _T_672; 
  wire [7:0] _T_673; 
  wire  _T_674; 
  wire  _T_675; 
  wire  _T_677; 
  wire  _T_678; 
  wire [7:0] _GEN_15; 
  wire  _T_682; 
  wire  _T_684; 
  wire  _T_685; 
  wire [7:0] _T_686; 
  wire [7:0] _T_687; 
  wire [7:0] _T_688; 
  wire  _T_689; 
  wire  _T_691; 
  wire  _T_692; 
  wire [7:0] _GEN_16; 
  wire  _T_693; 
  wire  _T_694; 
  wire  _T_695; 
  wire  _T_696; 
  wire  _T_698; 
  wire  _T_699; 
  wire [7:0] _T_700; 
  wire [7:0] _T_701; 
  wire [7:0] _T_702; 
  reg [31:0] _T_703; 
  reg [31:0] _RAND_16;
  wire  _T_704; 
  wire  _T_705; 
  wire  _T_706; 
  wire  _T_707; 
  wire  _T_708; 
  wire  _T_709; 
  wire  _T_711; 
  wire  _T_712; 
  wire [31:0] _T_714; 
  wire  _T_717; 
  wire  _GEN_19; 
  wire  _GEN_35; 
  wire  _GEN_53; 
  wire  _GEN_65; 
  wire  _GEN_75; 
  wire  _GEN_85; 
  wire  _GEN_95; 
  wire  _GEN_105; 
  wire  _GEN_115; 
  wire  _GEN_125; 
  wire  _GEN_137; 
  wire  _GEN_149; 
  wire  _GEN_155; 
  wire  _GEN_161; 
  dual_plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0)) plusarg_reader ( 
    .out(plusarg_reader_out)
  );
  assign _T_7 = io_in_a_bits_source[2:2]; 
  assign _T_8 = _T_7 == 1'h0; 
  assign _T_22 = _T_8 | _T_7; 
  assign _T_24 = 27'hfff << io_in_a_bits_size; 
  assign _T_25 = _T_24[11:0]; 
  assign _T_26 = ~ _T_25; 
  assign _GEN_18 = {{116'd0}, _T_26}; 
  assign _T_27 = io_in_a_bits_address & _GEN_18; 
  assign _T_28 = _T_27 == 128'h0; 
  assign _T_30 = io_in_a_bits_size[0]; 
  assign _T_31 = 2'h1 << _T_30; 
  assign _T_33 = _T_31 | 2'h1; 
  assign _T_34 = io_in_a_bits_size >= 4'h2; 
  assign _T_35 = _T_33[1]; 
  assign _T_36 = io_in_a_bits_address[1]; 
  assign _T_37 = _T_36 == 1'h0; 
  assign _T_39 = _T_35 & _T_37; 
  assign _T_40 = _T_34 | _T_39; 
  assign _T_42 = _T_35 & _T_36; 
  assign _T_43 = _T_34 | _T_42; 
  assign _T_44 = _T_33[0]; 
  assign _T_45 = io_in_a_bits_address[0]; 
  assign _T_46 = _T_45 == 1'h0; 
  assign _T_47 = _T_37 & _T_46; 
  assign _T_48 = _T_44 & _T_47; 
  assign _T_49 = _T_40 | _T_48; 
  assign _T_50 = _T_37 & _T_45; 
  assign _T_51 = _T_44 & _T_50; 
  assign _T_52 = _T_40 | _T_51; 
  assign _T_53 = _T_36 & _T_46; 
  assign _T_54 = _T_44 & _T_53; 
  assign _T_55 = _T_43 | _T_54; 
  assign _T_56 = _T_36 & _T_45; 
  assign _T_57 = _T_44 & _T_56; 
  assign _T_58 = _T_43 | _T_57; 
  assign _T_61 = {_T_58,_T_55,_T_52,_T_49}; 
  assign _T_72 = {1'b0,$signed(io_in_a_bits_address)}; 
  assign _T_96 = io_in_a_bits_opcode == 3'h6; 
  assign _T_98 = io_in_a_bits_size <= 4'hc; 
  assign _T_103 = $signed(_T_72) & $signed(-129'sh100000000000000000000000000000000); 
  assign _T_104 = $signed(_T_103); 
  assign _T_105 = $signed(_T_104) == $signed(129'sh0); 
  assign _T_106 = _T_98 & _T_105; 
  assign _T_109 = _T_106 | reset; 
  assign _T_110 = _T_109 == 1'h0; 
  assign _T_113 = reset == 1'h0; 
  assign _T_115 = _T_22 | reset; 
  assign _T_116 = _T_115 == 1'h0; 
  assign _T_119 = _T_34 | reset; 
  assign _T_120 = _T_119 == 1'h0; 
  assign _T_122 = _T_28 | reset; 
  assign _T_123 = _T_122 == 1'h0; 
  assign _T_124 = io_in_a_bits_param <= 3'h2; 
  assign _T_126 = _T_124 | reset; 
  assign _T_127 = _T_126 == 1'h0; 
  assign _T_128 = ~ io_in_a_bits_mask; 
  assign _T_129 = _T_128 == 4'h0; 
  assign _T_131 = _T_129 | reset; 
  assign _T_132 = _T_131 == 1'h0; 
  assign _T_133 = io_in_a_bits_corrupt == 1'h0; 
  assign _T_135 = _T_133 | reset; 
  assign _T_136 = _T_135 == 1'h0; 
  assign _T_137 = io_in_a_bits_opcode == 3'h7; 
  assign _T_169 = io_in_a_bits_param != 3'h0; 
  assign _T_171 = _T_169 | reset; 
  assign _T_172 = _T_171 == 1'h0; 
  assign _T_182 = io_in_a_bits_opcode == 3'h4; 
  assign _T_203 = io_in_a_bits_param == 3'h0; 
  assign _T_205 = _T_203 | reset; 
  assign _T_206 = _T_205 == 1'h0; 
  assign _T_207 = io_in_a_bits_mask == _T_61; 
  assign _T_209 = _T_207 | reset; 
  assign _T_210 = _T_209 == 1'h0; 
  assign _T_215 = io_in_a_bits_opcode == 3'h0; 
  assign _T_244 = io_in_a_bits_opcode == 3'h1; 
  assign _T_269 = ~ _T_61; 
  assign _T_270 = io_in_a_bits_mask & _T_269; 
  assign _T_271 = _T_270 == 4'h0; 
  assign _T_273 = _T_271 | reset; 
  assign _T_274 = _T_273 == 1'h0; 
  assign _T_275 = io_in_a_bits_opcode == 3'h2; 
  assign _T_277 = io_in_a_bits_size <= 4'h4; 
  assign _T_285 = _T_277 & _T_105; 
  assign _T_288 = _T_285 | reset; 
  assign _T_289 = _T_288 == 1'h0; 
  assign _T_296 = io_in_a_bits_param <= 3'h4; 
  assign _T_298 = _T_296 | reset; 
  assign _T_299 = _T_298 == 1'h0; 
  assign _T_304 = io_in_a_bits_opcode == 3'h3; 
  assign _T_325 = io_in_a_bits_param <= 3'h3; 
  assign _T_327 = _T_325 | reset; 
  assign _T_328 = _T_327 == 1'h0; 
  assign _T_333 = io_in_a_bits_opcode == 3'h5; 
  assign _T_362 = io_in_d_bits_opcode <= 3'h6; 
  assign _T_364 = _T_362 | reset; 
  assign _T_365 = _T_364 == 1'h0; 
  assign _T_368 = io_in_d_bits_source[2:2]; 
  assign _T_369 = _T_368 == 1'h0; 
  assign _T_383 = _T_369 | _T_368; 
  assign _T_384 = io_in_d_bits_sink < 1'h1; 
  assign _T_385 = io_in_d_bits_opcode == 3'h6; 
  assign _T_387 = _T_383 | reset; 
  assign _T_388 = _T_387 == 1'h0; 
  assign _T_389 = io_in_d_bits_size >= 4'h2; 
  assign _T_391 = _T_389 | reset; 
  assign _T_392 = _T_391 == 1'h0; 
  assign _T_393 = io_in_d_bits_param == 2'h0; 
  assign _T_395 = _T_393 | reset; 
  assign _T_396 = _T_395 == 1'h0; 
  assign _T_397 = io_in_d_bits_corrupt == 1'h0; 
  assign _T_399 = _T_397 | reset; 
  assign _T_400 = _T_399 == 1'h0; 
  assign _T_401 = io_in_d_bits_denied == 1'h0; 
  assign _T_403 = _T_401 | reset; 
  assign _T_404 = _T_403 == 1'h0; 
  assign _T_405 = io_in_d_bits_opcode == 3'h4; 
  assign _T_410 = _T_384 | reset; 
  assign _T_411 = _T_410 == 1'h0; 
  assign _T_416 = io_in_d_bits_param <= 2'h2; 
  assign _T_418 = _T_416 | reset; 
  assign _T_419 = _T_418 == 1'h0; 
  assign _T_420 = io_in_d_bits_param != 2'h2; 
  assign _T_422 = _T_420 | reset; 
  assign _T_423 = _T_422 == 1'h0; 
  assign _T_433 = io_in_d_bits_opcode == 3'h5; 
  assign _T_453 = _T_401 | io_in_d_bits_corrupt; 
  assign _T_455 = _T_453 | reset; 
  assign _T_456 = _T_455 == 1'h0; 
  assign _T_462 = io_in_d_bits_opcode == 3'h0; 
  assign _T_479 = io_in_d_bits_opcode == 3'h1; 
  assign _T_497 = io_in_d_bits_opcode == 3'h2; 
  assign _T_526 = io_in_a_ready & io_in_a_valid; 
  assign _T_531 = _T_26[11:2]; 
  assign _T_532 = io_in_a_bits_opcode[2]; 
  assign _T_533 = _T_532 == 1'h0; 
  assign _T_537 = _T_535 - 10'h1; 
  assign _T_538 = _T_535 == 10'h0; 
  assign _T_551 = _T_538 == 1'h0; 
  assign _T_552 = io_in_a_valid & _T_551; 
  assign _T_553 = io_in_a_bits_opcode == _T_546; 
  assign _T_555 = _T_553 | reset; 
  assign _T_556 = _T_555 == 1'h0; 
  assign _T_557 = io_in_a_bits_param == _T_547; 
  assign _T_559 = _T_557 | reset; 
  assign _T_560 = _T_559 == 1'h0; 
  assign _T_561 = io_in_a_bits_size == _T_548; 
  assign _T_563 = _T_561 | reset; 
  assign _T_564 = _T_563 == 1'h0; 
  assign _T_565 = io_in_a_bits_source == _T_549; 
  assign _T_567 = _T_565 | reset; 
  assign _T_568 = _T_567 == 1'h0; 
  assign _T_569 = io_in_a_bits_address == _T_550; 
  assign _T_571 = _T_569 | reset; 
  assign _T_572 = _T_571 == 1'h0; 
  assign _T_574 = _T_526 & _T_538; 
  assign _T_575 = io_in_d_ready & io_in_d_valid; 
  assign _T_577 = 27'hfff << io_in_d_bits_size; 
  assign _T_578 = _T_577[11:0]; 
  assign _T_579 = ~ _T_578; 
  assign _T_580 = _T_579[11:2]; 
  assign _T_581 = io_in_d_bits_opcode[0]; 
  assign _T_585 = _T_583 - 10'h1; 
  assign _T_586 = _T_583 == 10'h0; 
  assign _T_600 = _T_586 == 1'h0; 
  assign _T_601 = io_in_d_valid & _T_600; 
  assign _T_602 = io_in_d_bits_opcode == _T_594; 
  assign _T_604 = _T_602 | reset; 
  assign _T_605 = _T_604 == 1'h0; 
  assign _T_606 = io_in_d_bits_param == _T_595; 
  assign _T_608 = _T_606 | reset; 
  assign _T_609 = _T_608 == 1'h0; 
  assign _T_610 = io_in_d_bits_size == _T_596; 
  assign _T_612 = _T_610 | reset; 
  assign _T_613 = _T_612 == 1'h0; 
  assign _T_614 = io_in_d_bits_source == _T_597; 
  assign _T_616 = _T_614 | reset; 
  assign _T_617 = _T_616 == 1'h0; 
  assign _T_618 = io_in_d_bits_sink == _T_598; 
  assign _T_620 = _T_618 | reset; 
  assign _T_621 = _T_620 == 1'h0; 
  assign _T_622 = io_in_d_bits_denied == _T_599; 
  assign _T_624 = _T_622 | reset; 
  assign _T_625 = _T_624 == 1'h0; 
  assign _T_627 = _T_575 & _T_586; 
  assign _T_640 = _T_638 - 10'h1; 
  assign _T_641 = _T_638 == 10'h0; 
  assign _T_659 = _T_657 - 10'h1; 
  assign _T_660 = _T_657 == 10'h0; 
  assign _T_670 = _T_526 & _T_641; 
  assign _T_672 = 8'h1 << io_in_a_bits_source; 
  assign _T_673 = _T_628 >> io_in_a_bits_source; 
  assign _T_674 = _T_673[0]; 
  assign _T_675 = _T_674 == 1'h0; 
  assign _T_677 = _T_675 | reset; 
  assign _T_678 = _T_677 == 1'h0; 
  assign _GEN_15 = _T_670 ? _T_672 : 8'h0; 
  assign _T_682 = _T_575 & _T_660; 
  assign _T_684 = _T_385 == 1'h0; 
  assign _T_685 = _T_682 & _T_684; 
  assign _T_686 = 8'h1 << io_in_d_bits_source; 
  assign _T_687 = _GEN_15 | _T_628; 
  assign _T_688 = _T_687 >> io_in_d_bits_source; 
  assign _T_689 = _T_688[0]; 
  assign _T_691 = _T_689 | reset; 
  assign _T_692 = _T_691 == 1'h0; 
  assign _GEN_16 = _T_685 ? _T_686 : 8'h0; 
  assign _T_693 = _GEN_15 != _GEN_16; 
  assign _T_694 = _GEN_15 != 8'h0; 
  assign _T_695 = _T_694 == 1'h0; 
  assign _T_696 = _T_693 | _T_695; 
  assign _T_698 = _T_696 | reset; 
  assign _T_699 = _T_698 == 1'h0; 
  assign _T_700 = _T_628 | _GEN_15; 
  assign _T_701 = ~ _GEN_16; 
  assign _T_702 = _T_700 & _T_701; 
  assign _T_704 = _T_628 != 8'h0; 
  assign _T_705 = _T_704 == 1'h0; 
  assign _T_706 = plusarg_reader_out == 32'h0; 
  assign _T_707 = _T_705 | _T_706; 
  assign _T_708 = _T_703 < plusarg_reader_out; 
  assign _T_709 = _T_707 | _T_708; 
  assign _T_711 = _T_709 | reset; 
  assign _T_712 = _T_711 == 1'h0; 
  assign _T_714 = _T_703 + 32'h1; 
  assign _T_717 = _T_526 | _T_575; 
  assign _GEN_19 = io_in_a_valid & _T_96; 
  assign _GEN_35 = io_in_a_valid & _T_137; 
  assign _GEN_53 = io_in_a_valid & _T_182; 
  assign _GEN_65 = io_in_a_valid & _T_215; 
  assign _GEN_75 = io_in_a_valid & _T_244; 
  assign _GEN_85 = io_in_a_valid & _T_275; 
  assign _GEN_95 = io_in_a_valid & _T_304; 
  assign _GEN_105 = io_in_a_valid & _T_333; 
  assign _GEN_115 = io_in_d_valid & _T_385; 
  assign _GEN_125 = io_in_d_valid & _T_405; 
  assign _GEN_137 = io_in_d_valid & _T_433; 
  assign _GEN_149 = io_in_d_valid & _T_462; 
  assign _GEN_155 = io_in_d_valid & _T_479; 
  assign _GEN_161 = io_in_d_valid & _T_497; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_535 = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_546 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_547 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_548 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_549 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {4{`RANDOM}};
  _T_550 = _RAND_5[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_583 = _RAND_6[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_594 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_595 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_596 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_597 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_598 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_599 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_628 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_638 = _RAND_14[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_657 = _RAND_15[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_703 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_535 <= 10'h0;
    end else begin
      if (_T_526) begin
        if (_T_538) begin
          if (_T_533) begin
            _T_535 <= _T_531;
          end else begin
            _T_535 <= 10'h0;
          end
        end else begin
          _T_535 <= _T_537;
        end
      end
    end
    if (_T_574) begin
      _T_546 <= io_in_a_bits_opcode;
    end
    if (_T_574) begin
      _T_547 <= io_in_a_bits_param;
    end
    if (_T_574) begin
      _T_548 <= io_in_a_bits_size;
    end
    if (_T_574) begin
      _T_549 <= io_in_a_bits_source;
    end
    if (_T_574) begin
      _T_550 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_583 <= 10'h0;
    end else begin
      if (_T_575) begin
        if (_T_586) begin
          if (_T_581) begin
            _T_583 <= _T_580;
          end else begin
            _T_583 <= 10'h0;
          end
        end else begin
          _T_583 <= _T_585;
        end
      end
    end
    if (_T_627) begin
      _T_594 <= io_in_d_bits_opcode;
    end
    if (_T_627) begin
      _T_595 <= io_in_d_bits_param;
    end
    if (_T_627) begin
      _T_596 <= io_in_d_bits_size;
    end
    if (_T_627) begin
      _T_597 <= io_in_d_bits_source;
    end
    if (_T_627) begin
      _T_598 <= io_in_d_bits_sink;
    end
    if (_T_627) begin
      _T_599 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_628 <= 8'h0;
    end else begin
      _T_628 <= _T_702;
    end
    if (reset) begin
      _T_638 <= 10'h0;
    end else begin
      if (_T_526) begin
        if (_T_641) begin
          if (_T_533) begin
            _T_638 <= _T_531;
          end else begin
            _T_638 <= 10'h0;
          end
        end else begin
          _T_638 <= _T_640;
        end
      end
    end
    if (reset) begin
      _T_657 <= 10'h0;
    end else begin
      if (_T_575) begin
        if (_T_660) begin
          if (_T_581) begin
            _T_657 <= _T_580;
          end else begin
            _T_657 <= 10'h0;
          end
        end else begin
          _T_657 <= _T_659;
        end
      end
    end
    if (reset) begin
      _T_703 <= 32'h0;
    end else begin
      if (_T_717) begin
        _T_703 <= 32'h0;
      end else begin
        _T_703 <= _T_714;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel has invalid opcode (connected at BusBypass.scala:32:14)\n    at Monitor.scala:39 assert (TLMessages.isA(bundle.opcode), \"'A' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:46 assert (visible(edge.address(bundle), bundle.source, edge), \"'A' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at BusBypass.scala:32:14)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_110) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_113) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at BusBypass.scala:32:14)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_113) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at BusBypass.scala:32:14)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_120) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at BusBypass.scala:32:14)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_120) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_123) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at BusBypass.scala:32:14)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_123) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_127) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at BusBypass.scala:32:14)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_127) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_132) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at BusBypass.scala:32:14)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_132) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_136) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at BusBypass.scala:32:14)\n    at Monitor.scala:56 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_136) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at BusBypass.scala:32:14)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_110) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_113) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at BusBypass.scala:32:14)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_113) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at BusBypass.scala:32:14)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_120) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at BusBypass.scala:32:14)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_120) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_123) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at BusBypass.scala:32:14)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_123) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_127) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at BusBypass.scala:32:14)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_127) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_172) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at BusBypass.scala:32:14)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_172) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_132) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at BusBypass.scala:32:14)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_132) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_136) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at BusBypass.scala:32:14)\n    at Monitor.scala:68 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_136) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at BusBypass.scala:32:14)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_110) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at BusBypass.scala:32:14)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_123) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at BusBypass.scala:32:14)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_123) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_206) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at BusBypass.scala:32:14)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_206) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_210) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at BusBypass.scala:32:14)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_210) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_136) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at BusBypass.scala:32:14)\n    at Monitor.scala:77 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_136) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at BusBypass.scala:32:14)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_110) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at BusBypass.scala:32:14)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_123) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at BusBypass.scala:32:14)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_123) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_206) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at BusBypass.scala:32:14)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_206) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_210) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at BusBypass.scala:32:14)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_210) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at BusBypass.scala:32:14)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_110) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at BusBypass.scala:32:14)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_123) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at BusBypass.scala:32:14)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_123) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_206) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at BusBypass.scala:32:14)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_206) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_274) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at BusBypass.scala:32:14)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_274) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_289) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at BusBypass.scala:32:14)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_289) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at BusBypass.scala:32:14)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_123) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at BusBypass.scala:32:14)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_123) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_299) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at BusBypass.scala:32:14)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_299) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_210) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at BusBypass.scala:32:14)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_210) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_289) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at BusBypass.scala:32:14)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_289) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at BusBypass.scala:32:14)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_123) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at BusBypass.scala:32:14)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_123) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_328) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at BusBypass.scala:32:14)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_328) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_210) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at BusBypass.scala:32:14)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_210) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_110) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at BusBypass.scala:32:14)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_110) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at BusBypass.scala:32:14)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_123) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at BusBypass.scala:32:14)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_123) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_210) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at BusBypass.scala:32:14)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_210) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_136) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at BusBypass.scala:32:14)\n    at Monitor.scala:117 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_136) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_365) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at BusBypass.scala:32:14)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_365) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_388) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at BusBypass.scala:32:14)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_388) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_392) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at BusBypass.scala:32:14)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_392) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_396) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at BusBypass.scala:32:14)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_396) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_400) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at BusBypass.scala:32:14)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_400) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_404) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at BusBypass.scala:32:14)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_404) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_388) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at BusBypass.scala:32:14)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_388) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_411) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at BusBypass.scala:32:14)\n    at Monitor.scala:285 assert (sink_ok, \"'D' channel Grant carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_411) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_392) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at BusBypass.scala:32:14)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_392) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_419) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at BusBypass.scala:32:14)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_419) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_423) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at BusBypass.scala:32:14)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_423) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_400) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at BusBypass.scala:32:14)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_400) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is denied (connected at BusBypass.scala:32:14)\n    at Monitor.scala:290 assert (deny_put_ok || !bundle.denied, \"'D' channel Grant is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_388) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at BusBypass.scala:32:14)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_388) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_411) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at BusBypass.scala:32:14)\n    at Monitor.scala:295 assert (sink_ok, \"'D' channel GrantData carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_411) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_392) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at BusBypass.scala:32:14)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_392) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_419) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at BusBypass.scala:32:14)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_419) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_423) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at BusBypass.scala:32:14)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_423) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_456) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at BusBypass.scala:32:14)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_456) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied (connected at BusBypass.scala:32:14)\n    at Monitor.scala:300 assert (deny_get_ok || !bundle.denied, \"'D' channel GrantData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_388) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at BusBypass.scala:32:14)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_388) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_396) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at BusBypass.scala:32:14)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_396) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_400) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at BusBypass.scala:32:14)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_400) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is denied (connected at BusBypass.scala:32:14)\n    at Monitor.scala:308 assert (deny_put_ok || !bundle.denied, \"'D' channel AccessAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_388) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at BusBypass.scala:32:14)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_388) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_396) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at BusBypass.scala:32:14)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_396) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_456) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at BusBypass.scala:32:14)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_456) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied (connected at BusBypass.scala:32:14)\n    at Monitor.scala:316 assert (deny_get_ok || !bundle.denied, \"'D' channel AccessAckData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_388) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at BusBypass.scala:32:14)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_388) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_396) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at BusBypass.scala:32:14)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_396) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_400) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at BusBypass.scala:32:14)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_400) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is denied (connected at BusBypass.scala:32:14)\n    at Monitor.scala:324 assert (deny_put_ok || !bundle.denied, \"'D' channel HintAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel valid and not TL-C (connected at BusBypass.scala:32:14)\n    at Monitor.scala:341 assert (!bundle.b.valid, \"'B' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel valid and not TL-C (connected at BusBypass.scala:32:14)\n    at Monitor.scala:342 assert (!bundle.c.valid, \"'C' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel valid and not TL-C (connected at BusBypass.scala:32:14)\n    at Monitor.scala:343 assert (!bundle.e.valid, \"'E' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_552 & _T_556) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at BusBypass.scala:32:14)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_552 & _T_556) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_552 & _T_560) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at BusBypass.scala:32:14)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_552 & _T_560) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_552 & _T_564) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at BusBypass.scala:32:14)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_552 & _T_564) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_552 & _T_568) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at BusBypass.scala:32:14)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_552 & _T_568) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_552 & _T_572) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at BusBypass.scala:32:14)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_552 & _T_572) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_601 & _T_605) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at BusBypass.scala:32:14)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_601 & _T_605) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_601 & _T_609) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at BusBypass.scala:32:14)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_601 & _T_609) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_601 & _T_613) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at BusBypass.scala:32:14)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_601 & _T_613) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_601 & _T_617) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at BusBypass.scala:32:14)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_601 & _T_617) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_601 & _T_621) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at BusBypass.scala:32:14)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_601 & _T_621) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_601 & _T_625) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at BusBypass.scala:32:14)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_601 & _T_625) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_670 & _T_678) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at BusBypass.scala:32:14)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_670 & _T_678) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_685 & _T_692) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at BusBypass.scala:32:14)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_685 & _T_692) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_699) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at BusBypass.scala:32:14)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_699) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_712) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at BusBypass.scala:32:14)\n    at Monitor.scala:479 assert (!inflight.orR || limit === UInt(0) || watchdog < limit, \"TileLink timeout expired\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_712) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLMonitor_5( 
  input         clock, 
  input         reset, 
  input         io_in_c_ready, 
  input         io_in_c_valid, 
  input  [2:0]  io_in_c_bits_opcode, 
  input  [2:0]  io_in_c_bits_param, 
  input  [3:0]  io_in_c_bits_size, 
  input         io_in_c_bits_source, 
  input  [31:0] io_in_c_bits_address, 
  input         io_in_c_bits_corrupt, 
  input         io_in_d_valid, 
  input  [2:0]  io_in_d_bits_opcode, 
  input  [1:0]  io_in_d_bits_param, 
  input  [3:0]  io_in_d_bits_size, 
  input         io_in_d_bits_source, 
  input         io_in_d_bits_sink, 
  input         io_in_d_bits_denied, 
  input         io_in_d_bits_corrupt 
);
  wire [31:0] plusarg_reader_out; 
  wire  _T_444; 
  wire  _T_446; 
  wire  _T_447; 
  wire  _T_448; 
  wire  _T_450; 
  wire  _T_451; 
  wire  _T_453; 
  wire  _T_454; 
  wire  _T_455; 
  wire  _T_457; 
  wire  _T_458; 
  wire  _T_459; 
  wire  _T_461; 
  wire  _T_462; 
  wire  _T_463; 
  wire  _T_465; 
  wire  _T_466; 
  wire  _T_467; 
  wire  _T_469; 
  wire  _T_470; 
  wire  _T_471; 
  wire  _T_476; 
  wire  _T_477; 
  wire  _T_482; 
  wire  _T_484; 
  wire  _T_485; 
  wire  _T_486; 
  wire  _T_488; 
  wire  _T_489; 
  wire  _T_499; 
  wire  _T_519; 
  wire  _T_521; 
  wire  _T_522; 
  wire  _T_528; 
  wire  _T_545; 
  wire  _T_563; 
  wire  _T_819; 
  wire [22:0] _T_822; 
  wire [7:0] _T_823; 
  wire [7:0] _T_824; 
  wire [31:0] _GEN_33; 
  wire [31:0] _T_825; 
  wire  _T_826; 
  wire [31:0] _T_827; 
  wire [32:0] _T_828; 
  wire [32:0] _T_829; 
  wire [32:0] _T_830; 
  wire  _T_831; 
  wire [31:0] _T_832; 
  wire [32:0] _T_833; 
  wire [32:0] _T_834; 
  wire [32:0] _T_835; 
  wire  _T_836; 
  wire [31:0] _T_837; 
  wire [32:0] _T_838; 
  wire [32:0] _T_839; 
  wire [32:0] _T_840; 
  wire  _T_841; 
  wire  _T_843; 
  wire  _T_844; 
  wire  _T_856; 
  wire  _T_858; 
  wire  _T_859; 
  wire  _T_861; 
  wire  _T_862; 
  wire  _T_863; 
  wire  _T_865; 
  wire  _T_866; 
  wire  _T_868; 
  wire  _T_869; 
  wire  _T_870; 
  wire  _T_872; 
  wire  _T_873; 
  wire  _T_874; 
  wire  _T_876; 
  wire  _T_877; 
  wire  _T_878; 
  wire  _T_896; 
  wire  _T_911; 
  wire  _T_919; 
  wire  _T_923; 
  wire  _T_924; 
  wire  _T_929; 
  wire  _T_930; 
  wire  _T_941; 
  wire  _T_943; 
  wire  _T_944; 
  wire  _T_949; 
  wire  _T_998; 
  wire  _T_1008; 
  wire  _T_1010; 
  wire  _T_1011; 
  wire  _T_1016; 
  wire  _T_1030; 
  wire [22:0] _T_1103; 
  wire [7:0] _T_1104; 
  wire [7:0] _T_1105; 
  wire [5:0] _T_1106; 
  wire  _T_1107; 
  reg [5:0] _T_1109; 
  reg [31:0] _RAND_0;
  wire [5:0] _T_1111; 
  wire  _T_1112; 
  reg [2:0] _T_1120; 
  reg [31:0] _RAND_1;
  reg [1:0] _T_1121; 
  reg [31:0] _RAND_2;
  reg [3:0] _T_1122; 
  reg [31:0] _RAND_3;
  reg  _T_1123; 
  reg [31:0] _RAND_4;
  reg  _T_1124; 
  reg [31:0] _RAND_5;
  reg  _T_1125; 
  reg [31:0] _RAND_6;
  wire  _T_1126; 
  wire  _T_1127; 
  wire  _T_1128; 
  wire  _T_1130; 
  wire  _T_1131; 
  wire  _T_1132; 
  wire  _T_1134; 
  wire  _T_1135; 
  wire  _T_1136; 
  wire  _T_1138; 
  wire  _T_1139; 
  wire  _T_1140; 
  wire  _T_1142; 
  wire  _T_1143; 
  wire  _T_1144; 
  wire  _T_1146; 
  wire  _T_1147; 
  wire  _T_1148; 
  wire  _T_1150; 
  wire  _T_1151; 
  wire  _T_1153; 
  wire  _T_1203; 
  wire [5:0] _T_1208; 
  wire  _T_1209; 
  reg [5:0] _T_1211; 
  reg [31:0] _RAND_7;
  wire [5:0] _T_1213; 
  wire  _T_1214; 
  reg [2:0] _T_1222; 
  reg [31:0] _RAND_8;
  reg [2:0] _T_1223; 
  reg [31:0] _RAND_9;
  reg [3:0] _T_1224; 
  reg [31:0] _RAND_10;
  reg  _T_1225; 
  reg [31:0] _RAND_11;
  reg [31:0] _T_1226; 
  reg [31:0] _RAND_12;
  wire  _T_1227; 
  wire  _T_1228; 
  wire  _T_1229; 
  wire  _T_1231; 
  wire  _T_1232; 
  wire  _T_1233; 
  wire  _T_1235; 
  wire  _T_1236; 
  wire  _T_1237; 
  wire  _T_1239; 
  wire  _T_1240; 
  wire  _T_1241; 
  wire  _T_1243; 
  wire  _T_1244; 
  wire  _T_1245; 
  wire  _T_1247; 
  wire  _T_1248; 
  wire  _T_1250; 
  reg  _T_1251; 
  reg [31:0] _RAND_13;
  reg [5:0] _T_1280; 
  reg [31:0] _RAND_14;
  wire [5:0] _T_1282; 
  wire  _T_1283; 
  wire  _T_1298; 
  wire  _T_1305; 
  wire  _T_1307; 
  wire  _T_1308; 
  wire [1:0] _T_1309; 
  wire  _T_1311; 
  wire  _T_1314; 
  wire  _T_1315; 
  wire [1:0] _GEN_28; 
  wire  _T_1302; 
  wire  _T_1324; 
  wire  _T_1325; 
  reg [31:0] _T_1326; 
  reg [31:0] _RAND_15;
  wire  _T_1329; 
  wire  _T_1330; 
  wire  _T_1331; 
  wire  _T_1332; 
  wire  _T_1334; 
  wire  _T_1335; 
  wire [31:0] _T_1337; 
  reg  _T_1341; 
  reg [31:0] _RAND_16;
  reg [5:0] _T_1350; 
  reg [31:0] _RAND_17;
  wire [5:0] _T_1352; 
  wire  _T_1353; 
  wire  _T_1363; 
  wire  _T_1364; 
  wire  _T_1365; 
  wire  _T_1366; 
  wire  _T_1367; 
  wire  _T_1368; 
  wire [1:0] _T_1369; 
  wire  _T_1370; 
  wire  _T_1372; 
  wire  _T_1374; 
  wire  _T_1375; 
  wire [1:0] _GEN_31; 
  wire  _T_1361; 
  wire  _T_1387; 
  wire  _GEN_34; 
  wire  _GEN_44; 
  wire  _GEN_56; 
  wire  _GEN_68; 
  wire  _GEN_74; 
  wire  _GEN_80; 
  wire  _GEN_86; 
  wire  _GEN_98; 
  wire  _GEN_108; 
  wire  _GEN_122; 
  wire  _GEN_134; 
  wire  _GEN_144; 
  wire  _GEN_152; 
  dual_plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0)) plusarg_reader ( 
    .out(plusarg_reader_out)
  );
  assign _T_444 = io_in_d_bits_opcode <= 3'h6; 
  assign _T_446 = _T_444 | reset; 
  assign _T_447 = _T_446 == 1'h0; 
  assign _T_448 = io_in_d_bits_source == 1'h0; 
  assign _T_450 = io_in_d_bits_sink < 1'h1; 
  assign _T_451 = io_in_d_bits_opcode == 3'h6; 
  assign _T_453 = _T_448 | reset; 
  assign _T_454 = _T_453 == 1'h0; 
  assign _T_455 = io_in_d_bits_size >= 4'h2; 
  assign _T_457 = _T_455 | reset; 
  assign _T_458 = _T_457 == 1'h0; 
  assign _T_459 = io_in_d_bits_param == 2'h0; 
  assign _T_461 = _T_459 | reset; 
  assign _T_462 = _T_461 == 1'h0; 
  assign _T_463 = io_in_d_bits_corrupt == 1'h0; 
  assign _T_465 = _T_463 | reset; 
  assign _T_466 = _T_465 == 1'h0; 
  assign _T_467 = io_in_d_bits_denied == 1'h0; 
  assign _T_469 = _T_467 | reset; 
  assign _T_470 = _T_469 == 1'h0; 
  assign _T_471 = io_in_d_bits_opcode == 3'h4; 
  assign _T_476 = _T_450 | reset; 
  assign _T_477 = _T_476 == 1'h0; 
  assign _T_482 = io_in_d_bits_param <= 2'h2; 
  assign _T_484 = _T_482 | reset; 
  assign _T_485 = _T_484 == 1'h0; 
  assign _T_486 = io_in_d_bits_param != 2'h2; 
  assign _T_488 = _T_486 | reset; 
  assign _T_489 = _T_488 == 1'h0; 
  assign _T_499 = io_in_d_bits_opcode == 3'h5; 
  assign _T_519 = _T_467 | io_in_d_bits_corrupt; 
  assign _T_521 = _T_519 | reset; 
  assign _T_522 = _T_521 == 1'h0; 
  assign _T_528 = io_in_d_bits_opcode == 3'h0; 
  assign _T_545 = io_in_d_bits_opcode == 3'h1; 
  assign _T_563 = io_in_d_bits_opcode == 3'h2; 
  assign _T_819 = io_in_c_bits_source == 1'h0; 
  assign _T_822 = 23'hff << io_in_c_bits_size; 
  assign _T_823 = _T_822[7:0]; 
  assign _T_824 = ~ _T_823; 
  assign _GEN_33 = {{24'd0}, _T_824}; 
  assign _T_825 = io_in_c_bits_address & _GEN_33; 
  assign _T_826 = _T_825 == 32'h0; 
  assign _T_827 = io_in_c_bits_address ^ 32'h80000000; 
  assign _T_828 = {1'b0,$signed(_T_827)}; 
  assign _T_829 = $signed(_T_828) & $signed(-33'sh80000000); 
  assign _T_830 = $signed(_T_829); 
  assign _T_831 = $signed(_T_830) == $signed(33'sh0); 
  assign _T_832 = io_in_c_bits_address ^ 32'h40000000; 
  assign _T_833 = {1'b0,$signed(_T_832)}; 
  assign _T_834 = $signed(_T_833) & $signed(-33'sh20000000); 
  assign _T_835 = $signed(_T_834); 
  assign _T_836 = $signed(_T_835) == $signed(33'sh0); 
  assign _T_837 = io_in_c_bits_address ^ 32'h10000000; 
  assign _T_838 = {1'b0,$signed(_T_837)}; 
  assign _T_839 = $signed(_T_838) & $signed(-33'sh10000000); 
  assign _T_840 = $signed(_T_839); 
  assign _T_841 = $signed(_T_840) == $signed(33'sh0); 
  assign _T_843 = _T_831 | _T_836; 
  assign _T_844 = _T_843 | _T_841; 
  assign _T_856 = io_in_c_bits_opcode == 3'h4; 
  assign _T_858 = _T_844 | reset; 
  assign _T_859 = _T_858 == 1'h0; 
  assign _T_861 = _T_819 | reset; 
  assign _T_862 = _T_861 == 1'h0; 
  assign _T_863 = io_in_c_bits_size >= 4'h2; 
  assign _T_865 = _T_863 | reset; 
  assign _T_866 = _T_865 == 1'h0; 
  assign _T_868 = _T_826 | reset; 
  assign _T_869 = _T_868 == 1'h0; 
  assign _T_870 = io_in_c_bits_param <= 3'h5; 
  assign _T_872 = _T_870 | reset; 
  assign _T_873 = _T_872 == 1'h0; 
  assign _T_874 = io_in_c_bits_corrupt == 1'h0; 
  assign _T_876 = _T_874 | reset; 
  assign _T_877 = _T_876 == 1'h0; 
  assign _T_878 = io_in_c_bits_opcode == 3'h5; 
  assign _T_896 = io_in_c_bits_opcode == 3'h6; 
  assign _T_911 = io_in_c_bits_size <= 4'h6; 
  assign _T_919 = _T_911 & _T_841; 
  assign _T_923 = _T_919 | reset; 
  assign _T_924 = _T_923 == 1'h0; 
  assign _T_929 = _T_911 | reset; 
  assign _T_930 = _T_929 == 1'h0; 
  assign _T_941 = io_in_c_bits_param <= 3'h2; 
  assign _T_943 = _T_941 | reset; 
  assign _T_944 = _T_943 == 1'h0; 
  assign _T_949 = io_in_c_bits_opcode == 3'h7; 
  assign _T_998 = io_in_c_bits_opcode == 3'h0; 
  assign _T_1008 = io_in_c_bits_param == 3'h0; 
  assign _T_1010 = _T_1008 | reset; 
  assign _T_1011 = _T_1010 == 1'h0; 
  assign _T_1016 = io_in_c_bits_opcode == 3'h1; 
  assign _T_1030 = io_in_c_bits_opcode == 3'h2; 
  assign _T_1103 = 23'hff << io_in_d_bits_size; 
  assign _T_1104 = _T_1103[7:0]; 
  assign _T_1105 = ~ _T_1104; 
  assign _T_1106 = _T_1105[7:2]; 
  assign _T_1107 = io_in_d_bits_opcode[0]; 
  assign _T_1111 = _T_1109 - 6'h1; 
  assign _T_1112 = _T_1109 == 6'h0; 
  assign _T_1126 = _T_1112 == 1'h0; 
  assign _T_1127 = io_in_d_valid & _T_1126; 
  assign _T_1128 = io_in_d_bits_opcode == _T_1120; 
  assign _T_1130 = _T_1128 | reset; 
  assign _T_1131 = _T_1130 == 1'h0; 
  assign _T_1132 = io_in_d_bits_param == _T_1121; 
  assign _T_1134 = _T_1132 | reset; 
  assign _T_1135 = _T_1134 == 1'h0; 
  assign _T_1136 = io_in_d_bits_size == _T_1122; 
  assign _T_1138 = _T_1136 | reset; 
  assign _T_1139 = _T_1138 == 1'h0; 
  assign _T_1140 = io_in_d_bits_source == _T_1123; 
  assign _T_1142 = _T_1140 | reset; 
  assign _T_1143 = _T_1142 == 1'h0; 
  assign _T_1144 = io_in_d_bits_sink == _T_1124; 
  assign _T_1146 = _T_1144 | reset; 
  assign _T_1147 = _T_1146 == 1'h0; 
  assign _T_1148 = io_in_d_bits_denied == _T_1125; 
  assign _T_1150 = _T_1148 | reset; 
  assign _T_1151 = _T_1150 == 1'h0; 
  assign _T_1153 = io_in_d_valid & _T_1112; 
  assign _T_1203 = io_in_c_ready & io_in_c_valid; 
  assign _T_1208 = _T_824[7:2]; 
  assign _T_1209 = io_in_c_bits_opcode[0]; 
  assign _T_1213 = _T_1211 - 6'h1; 
  assign _T_1214 = _T_1211 == 6'h0; 
  assign _T_1227 = _T_1214 == 1'h0; 
  assign _T_1228 = io_in_c_valid & _T_1227; 
  assign _T_1229 = io_in_c_bits_opcode == _T_1222; 
  assign _T_1231 = _T_1229 | reset; 
  assign _T_1232 = _T_1231 == 1'h0; 
  assign _T_1233 = io_in_c_bits_param == _T_1223; 
  assign _T_1235 = _T_1233 | reset; 
  assign _T_1236 = _T_1235 == 1'h0; 
  assign _T_1237 = io_in_c_bits_size == _T_1224; 
  assign _T_1239 = _T_1237 | reset; 
  assign _T_1240 = _T_1239 == 1'h0; 
  assign _T_1241 = io_in_c_bits_source == _T_1225; 
  assign _T_1243 = _T_1241 | reset; 
  assign _T_1244 = _T_1243 == 1'h0; 
  assign _T_1245 = io_in_c_bits_address == _T_1226; 
  assign _T_1247 = _T_1245 | reset; 
  assign _T_1248 = _T_1247 == 1'h0; 
  assign _T_1250 = _T_1203 & _T_1214; 
  assign _T_1282 = _T_1280 - 6'h1; 
  assign _T_1283 = _T_1280 == 6'h0; 
  assign _T_1298 = _T_1251 == 1'h0; 
  assign _T_1305 = io_in_d_valid & _T_1283; 
  assign _T_1307 = _T_451 == 1'h0; 
  assign _T_1308 = _T_1305 & _T_1307; 
  assign _T_1309 = 2'h1 << io_in_d_bits_source; 
  assign _T_1311 = _T_1251 >> io_in_d_bits_source; 
  assign _T_1314 = _T_1311 | reset; 
  assign _T_1315 = _T_1314 == 1'h0; 
  assign _GEN_28 = _T_1308 ? _T_1309 : 2'h0; 
  assign _T_1302 = _GEN_28[0]; 
  assign _T_1324 = ~ _T_1302; 
  assign _T_1325 = _T_1251 & _T_1324; 
  assign _T_1329 = plusarg_reader_out == 32'h0; 
  assign _T_1330 = _T_1298 | _T_1329; 
  assign _T_1331 = _T_1326 < plusarg_reader_out; 
  assign _T_1332 = _T_1330 | _T_1331; 
  assign _T_1334 = _T_1332 | reset; 
  assign _T_1335 = _T_1334 == 1'h0; 
  assign _T_1337 = _T_1326 + 32'h1; 
  assign _T_1352 = _T_1350 - 6'h1; 
  assign _T_1353 = _T_1350 == 6'h0; 
  assign _T_1363 = io_in_d_valid & _T_1353; 
  assign _T_1364 = io_in_d_bits_opcode[2]; 
  assign _T_1365 = io_in_d_bits_opcode[1]; 
  assign _T_1366 = _T_1365 == 1'h0; 
  assign _T_1367 = _T_1364 & _T_1366; 
  assign _T_1368 = _T_1363 & _T_1367; 
  assign _T_1369 = 2'h1 << io_in_d_bits_sink; 
  assign _T_1370 = _T_1341 >> io_in_d_bits_sink; 
  assign _T_1372 = _T_1370 == 1'h0; 
  assign _T_1374 = _T_1372 | reset; 
  assign _T_1375 = _T_1374 == 1'h0; 
  assign _GEN_31 = _T_1368 ? _T_1369 : 2'h0; 
  assign _T_1361 = _GEN_31[0]; 
  assign _T_1387 = _T_1341 | _T_1361; 
  assign _GEN_34 = io_in_d_valid & _T_451; 
  assign _GEN_44 = io_in_d_valid & _T_471; 
  assign _GEN_56 = io_in_d_valid & _T_499; 
  assign _GEN_68 = io_in_d_valid & _T_528; 
  assign _GEN_74 = io_in_d_valid & _T_545; 
  assign _GEN_80 = io_in_d_valid & _T_563; 
  assign _GEN_86 = io_in_c_valid & _T_856; 
  assign _GEN_98 = io_in_c_valid & _T_878; 
  assign _GEN_108 = io_in_c_valid & _T_896; 
  assign _GEN_122 = io_in_c_valid & _T_949; 
  assign _GEN_134 = io_in_c_valid & _T_998; 
  assign _GEN_144 = io_in_c_valid & _T_1016; 
  assign _GEN_152 = io_in_c_valid & _T_1030; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1109 = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1120 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1121 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1122 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1123 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1124 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_1125 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_1211 = _RAND_7[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1222 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_1223 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_1224 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_1225 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_1226 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_1251 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_1280 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_1326 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_1341 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_1350 = _RAND_17[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_1109 <= 6'h0;
    end else begin
      if (io_in_d_valid) begin
        if (_T_1112) begin
          if (_T_1107) begin
            _T_1109 <= _T_1106;
          end else begin
            _T_1109 <= 6'h0;
          end
        end else begin
          _T_1109 <= _T_1111;
        end
      end
    end
    if (_T_1153) begin
      _T_1120 <= io_in_d_bits_opcode;
    end
    if (_T_1153) begin
      _T_1121 <= io_in_d_bits_param;
    end
    if (_T_1153) begin
      _T_1122 <= io_in_d_bits_size;
    end
    if (_T_1153) begin
      _T_1123 <= io_in_d_bits_source;
    end
    if (_T_1153) begin
      _T_1124 <= io_in_d_bits_sink;
    end
    if (_T_1153) begin
      _T_1125 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_1211 <= 6'h0;
    end else begin
      if (_T_1203) begin
        if (_T_1214) begin
          if (_T_1209) begin
            _T_1211 <= _T_1208;
          end else begin
            _T_1211 <= 6'h0;
          end
        end else begin
          _T_1211 <= _T_1213;
        end
      end
    end
    if (_T_1250) begin
      _T_1222 <= io_in_c_bits_opcode;
    end
    if (_T_1250) begin
      _T_1223 <= io_in_c_bits_param;
    end
    if (_T_1250) begin
      _T_1224 <= io_in_c_bits_size;
    end
    if (_T_1250) begin
      _T_1225 <= io_in_c_bits_source;
    end
    if (_T_1250) begin
      _T_1226 <= io_in_c_bits_address;
    end
    if (reset) begin
      _T_1251 <= 1'h0;
    end else begin
      _T_1251 <= _T_1325;
    end
    if (reset) begin
      _T_1280 <= 6'h0;
    end else begin
      if (io_in_d_valid) begin
        if (_T_1283) begin
          if (_T_1107) begin
            _T_1280 <= _T_1106;
          end else begin
            _T_1280 <= 6'h0;
          end
        end else begin
          _T_1280 <= _T_1282;
        end
      end
    end
    if (reset) begin
      _T_1326 <= 32'h0;
    end else begin
      if (io_in_d_valid) begin
        _T_1326 <= 32'h0;
      end else begin
        _T_1326 <= _T_1337;
      end
    end
    if (reset) begin
      _T_1341 <= 1'h0;
    end else begin
      _T_1341 <= _T_1387;
    end
    if (reset) begin
      _T_1350 <= 6'h0;
    end else begin
      if (io_in_d_valid) begin
        if (_T_1353) begin
          if (_T_1107) begin
            _T_1350 <= _T_1106;
          end else begin
            _T_1350 <= 6'h0;
          end
        end else begin
          _T_1350 <= _T_1352;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel has invalid opcode (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:39 assert (TLMessages.isA(bundle.opcode), \"'A' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:46 assert (visible(edge.address(bundle), bundle.source, edge), \"'A' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:56 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:68 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:77 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:117 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_447) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_447) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_34 & _T_454) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_34 & _T_454) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_34 & _T_458) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_34 & _T_458) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_34 & _T_462) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_34 & _T_462) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_34 & _T_466) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_34 & _T_466) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_34 & _T_470) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_34 & _T_470) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_44 & _T_454) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_44 & _T_454) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_44 & _T_477) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:285 assert (sink_ok, \"'D' channel Grant carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_44 & _T_477) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_44 & _T_458) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_44 & _T_458) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_44 & _T_485) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_44 & _T_485) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_44 & _T_489) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_44 & _T_489) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_44 & _T_466) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_44 & _T_466) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is denied (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:290 assert (deny_put_ok || !bundle.denied, \"'D' channel Grant is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_454) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_56 & _T_454) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_477) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:295 assert (sink_ok, \"'D' channel GrantData carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_56 & _T_477) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_458) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_56 & _T_458) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_485) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_56 & _T_485) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_489) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_56 & _T_489) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_522) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_56 & _T_522) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:300 assert (deny_get_ok || !bundle.denied, \"'D' channel GrantData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_68 & _T_454) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_68 & _T_454) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_68 & _T_462) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_68 & _T_462) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_68 & _T_466) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_68 & _T_466) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is denied (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:308 assert (deny_put_ok || !bundle.denied, \"'D' channel AccessAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_74 & _T_454) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_74 & _T_454) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_74 & _T_462) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_74 & _T_462) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_74 & _T_522) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_74 & _T_522) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:316 assert (deny_get_ok || !bundle.denied, \"'D' channel AccessAckData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_80 & _T_454) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_80 & _T_454) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_80 & _T_462) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_80 & _T_462) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_80 & _T_466) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_80 & _T_466) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is denied (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:324 assert (deny_put_ok || !bundle.denied, \"'D' channel HintAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel has invalid opcode (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:122 assert (TLMessages.isB(bundle.opcode), \"'B' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:124 assert (visible(edge.address(bundle), bundle.source, edge), \"'B' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Probe type unsupported by client (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:133 assert (edge.client.supportsProbe(bundle.source, bundle.size), \"'B' channel carries Probe type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:134 assert (address_ok, \"'B' channel Probe carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries source that is not first source (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:135 assert (legal_source, \"'B' channel Probe carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:136 assert (is_aligned, \"'B' channel Probe address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:137 assert (TLPermissions.isCap(bundle.param), \"'B' channel Probe carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe contains invalid mask (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:138 assert (bundle.mask === mask, \"'B' channel Probe contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe is corrupt (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:139 assert (!bundle.corrupt, \"'B' channel Probe is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Get type unsupported by client (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:143 assert (edge.client.supportsGet(bundle.source, bundle.size), \"'B' channel carries Get type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries unmanaged address (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:144 assert (address_ok, \"'B' channel Get carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries source that is not first source (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:145 assert (legal_source, \"'B' channel Get carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:146 assert (is_aligned, \"'B' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries invalid param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:147 assert (bundle.param === UInt(0), \"'B' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get contains invalid mask (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:148 assert (bundle.mask === mask, \"'B' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get is corrupt (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:149 assert (!bundle.corrupt, \"'B' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutFull type unsupported by client (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:153 assert (edge.client.supportsPutFull(bundle.source, bundle.size), \"'B' channel carries PutFull type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries unmanaged address (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:154 assert (address_ok, \"'B' channel PutFull carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries source that is not first source (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:155 assert (legal_source, \"'B' channel PutFull carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:156 assert (is_aligned, \"'B' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries invalid param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:157 assert (bundle.param === UInt(0), \"'B' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull contains invalid mask (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:158 assert (bundle.mask === mask, \"'B' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutPartial type unsupported by client (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:162 assert (edge.client.supportsPutPartial(bundle.source, bundle.size), \"'B' channel carries PutPartial type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:163 assert (address_ok, \"'B' channel PutPartial carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:164 assert (legal_source, \"'B' channel PutPartial carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:165 assert (is_aligned, \"'B' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries invalid param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:166 assert (bundle.param === UInt(0), \"'B' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial contains invalid mask (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:167 assert ((bundle.mask & ~mask) === UInt(0), \"'B' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Arithmetic type unsupported by client (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:171 assert (edge.client.supportsArithmetic(bundle.source, bundle.size), \"'B' channel carries Arithmetic type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:172 assert (address_ok, \"'B' channel Arithmetic carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:173 assert (legal_source, \"'B' channel Arithmetic carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:174 assert (is_aligned, \"'B' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries invalid opcode param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:175 assert (TLAtomics.isArithmetic(bundle.param), \"'B' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:176 assert (bundle.mask === mask, \"'B' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Logical type unsupported by client (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:180 assert (edge.client.supportsLogical(bundle.source, bundle.size), \"'B' channel carries Logical type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries unmanaged address (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:181 assert (address_ok, \"'B' channel Logical carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries source that is not first source (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:182 assert (legal_source, \"'B' channel Logical carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:183 assert (is_aligned, \"'B' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries invalid opcode param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:184 assert (TLAtomics.isLogical(bundle.param), \"'B' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical contains invalid mask (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:185 assert (bundle.mask === mask, \"'B' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Hint type unsupported by client (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:189 assert (edge.client.supportsHint(bundle.source, bundle.size), \"'B' channel carries Hint type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries unmanaged address (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:190 assert (address_ok, \"'B' channel Hint carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries source that is not first source (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:191 assert (legal_source, \"'B' channel Hint carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:192 assert (is_aligned, \"'B' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint contains invalid mask (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:193 assert (bundle.mask === mask, \"'B' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint is corrupt (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:194 assert (!bundle.corrupt, \"'B' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel has invalid opcode (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:199 assert (TLMessages.isC(bundle.opcode), \"'C' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:205 assert (visible(edge.address(bundle), bundle.source, edge), \"'C' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_86 & _T_859) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:208 assert (address_ok, \"'C' channel ProbeAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_86 & _T_859) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_86 & _T_862) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:209 assert (source_ok, \"'C' channel ProbeAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_86 & _T_862) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_86 & _T_866) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:210 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_86 & _T_866) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_86 & _T_869) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:211 assert (is_aligned, \"'C' channel ProbeAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_86 & _T_869) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_86 & _T_873) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:212 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAck carries invalid report param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_86 & _T_873) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_86 & _T_877) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck is corrupt (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:213 assert (!bundle.corrupt, \"'C' channel ProbeAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_86 & _T_877) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_859) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:217 assert (address_ok, \"'C' channel ProbeAckData carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_859) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_862) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:218 assert (source_ok, \"'C' channel ProbeAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_862) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_866) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:219 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAckData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_866) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_869) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:220 assert (is_aligned, \"'C' channel ProbeAckData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_869) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_873) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:221 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAckData carries invalid report param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_873) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_108 & _T_924) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:225 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries Release type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_108 & _T_924) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_108 & _T_930) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:226 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_108 & _T_930) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_108 & _T_862) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:227 assert (source_ok, \"'C' channel Release carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_108 & _T_862) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_108 & _T_866) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:228 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel Release smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_108 & _T_866) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_108 & _T_869) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:229 assert (is_aligned, \"'C' channel Release address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_108 & _T_869) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_108 & _T_944) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid shrink param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:230 assert (TLPermissions.isShrink(bundle.param), \"'C' channel Release carries invalid shrink param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_108 & _T_944) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_108 & _T_877) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release is corrupt (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:231 assert (!bundle.corrupt, \"'C' channel Release is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_108 & _T_877) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_122 & _T_924) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:235 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries ReleaseData type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_122 & _T_924) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_122 & _T_930) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:236 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_122 & _T_930) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_122 & _T_862) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:237 assert (source_ok, \"'C' channel ReleaseData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_122 & _T_862) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_122 & _T_866) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:238 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ReleaseData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_122 & _T_866) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_122 & _T_869) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:239 assert (is_aligned, \"'C' channel ReleaseData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_122 & _T_869) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_122 & _T_944) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid shrink param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:240 assert (TLPermissions.isShrink(bundle.param), \"'C' channel ReleaseData carries invalid shrink param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_122 & _T_944) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_134 & _T_859) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:244 assert (address_ok, \"'C' channel AccessAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_134 & _T_859) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_134 & _T_862) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:245 assert (source_ok, \"'C' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_134 & _T_862) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_134 & _T_869) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:246 assert (is_aligned, \"'C' channel AccessAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_134 & _T_869) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_134 & _T_1011) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:247 assert (bundle.param === UInt(0), \"'C' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_134 & _T_1011) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_134 & _T_877) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck is corrupt (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:248 assert (!bundle.corrupt, \"'C' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_134 & _T_877) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & _T_859) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:252 assert (address_ok, \"'C' channel AccessAckData carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_859) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & _T_862) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:253 assert (source_ok, \"'C' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_862) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & _T_869) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:254 assert (is_aligned, \"'C' channel AccessAckData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_869) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & _T_1011) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:255 assert (bundle.param === UInt(0), \"'C' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_1011) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_152 & _T_859) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:259 assert (address_ok, \"'C' channel HintAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_152 & _T_859) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_152 & _T_862) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:260 assert (source_ok, \"'C' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_152 & _T_862) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_152 & _T_869) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:261 assert (is_aligned, \"'C' channel HintAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_152 & _T_869) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_152 & _T_1011) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:262 assert (bundle.param === UInt(0), \"'C' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_152 & _T_1011) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_152 & _T_877) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck is corrupt (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:263 assert (!bundle.corrupt, \"'C' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_152 & _T_877) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channels carries invalid sink ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:330 assert (sink_ok, \"'E' channels carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1127 & _T_1131) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1127 & _T_1131) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1127 & _T_1135) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1127 & _T_1135) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1127 & _T_1139) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1127 & _T_1139) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1127 & _T_1143) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1127 & _T_1143) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1127 & _T_1147) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1127 & _T_1147) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1127 & _T_1151) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1127 & _T_1151) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel opcode changed within multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:378 assert (b.bits.opcode === opcode, \"'B' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:379 assert (b.bits.param  === param,  \"'B' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel size changed within multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:380 assert (b.bits.size   === size,   \"'B' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel source changed within multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:381 assert (b.bits.source === source, \"'B' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:382 assert (b.bits.address=== address,\"'B' channel addresss changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1228 & _T_1232) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:401 assert (c.bits.opcode === opcode, \"'C' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1228 & _T_1232) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1228 & _T_1236) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:402 assert (c.bits.param  === param,  \"'C' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1228 & _T_1236) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1228 & _T_1240) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:403 assert (c.bits.size   === size,   \"'C' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1228 & _T_1240) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1228 & _T_1244) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:404 assert (c.bits.source === source, \"'C' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1228 & _T_1244) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1228 & _T_1248) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:405 assert (c.bits.address=== address,\"'C' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1228 & _T_1248) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1308 & _T_1315) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1308 & _T_1315) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1335) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:479 assert (!inflight.orR || limit === UInt(0) || watchdog < limit, \"TileLink timeout expired\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1335) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1368 & _T_1375) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:494 assert(!inflight(bundle.d.bits.sink), \"'D' channel re-used a sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1368 & _T_1375) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at dual_ChipLink.scala:77:16)\n    at Monitor.scala:500 assert((d_set | inflight)(bundle.e.bits.sink), \"'E' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLMonitor_6( 
  input         clock, 
  input         reset, 
  input         io_in_a_ready, 
  input         io_in_a_valid, 
  input  [2:0]  io_in_a_bits_opcode, 
  input  [2:0]  io_in_a_bits_param, 
  input  [3:0]  io_in_a_bits_size, 
  input  [5:0]  io_in_a_bits_source, 
  input  [31:0] io_in_a_bits_address, 
  input  [3:0]  io_in_a_bits_mask, 
  input         io_in_c_ready, 
  input         io_in_c_valid, 
  input  [2:0]  io_in_c_bits_opcode, 
  input  [2:0]  io_in_c_bits_param, 
  input  [3:0]  io_in_c_bits_size, 
  input  [5:0]  io_in_c_bits_source, 
  input  [31:0] io_in_c_bits_address, 
  input         io_in_d_ready, 
  input         io_in_d_valid, 
  input  [2:0]  io_in_d_bits_opcode, 
  input  [1:0]  io_in_d_bits_param, 
  input  [3:0]  io_in_d_bits_size, 
  input  [5:0]  io_in_d_bits_source, 
  input         io_in_d_bits_sink, 
  input         io_in_d_bits_denied, 
  input         io_in_d_bits_corrupt, 
  input         io_in_e_ready, 
  input         io_in_e_valid, 
  input         io_in_e_bits_sink 
);
  wire [31:0] plusarg_reader_out; 
  wire [2:0] _T_7; 
  wire  _T_8; 
  wire  _T_16; 
  wire  _T_24; 
  wire  _T_32; 
  wire  _T_40; 
  wire  _T_48; 
  wire  _T_56; 
  wire  _T_64; 
  wire  _T_70; 
  wire  _T_71; 
  wire  _T_72; 
  wire  _T_73; 
  wire  _T_74; 
  wire  _T_75; 
  wire  _T_76; 
  wire [22:0] _T_78; 
  wire [7:0] _T_79; 
  wire [7:0] _T_80; 
  wire [31:0] _GEN_33; 
  wire [31:0] _T_81; 
  wire  _T_82; 
  wire  _T_84; 
  wire [1:0] _T_85; 
  wire [1:0] _T_87; 
  wire  _T_88; 
  wire  _T_89; 
  wire  _T_90; 
  wire  _T_91; 
  wire  _T_93; 
  wire  _T_94; 
  wire  _T_96; 
  wire  _T_97; 
  wire  _T_98; 
  wire  _T_99; 
  wire  _T_100; 
  wire  _T_101; 
  wire  _T_102; 
  wire  _T_103; 
  wire  _T_104; 
  wire  _T_105; 
  wire  _T_106; 
  wire  _T_107; 
  wire  _T_108; 
  wire  _T_109; 
  wire  _T_110; 
  wire  _T_111; 
  wire  _T_112; 
  wire [3:0] _T_115; 
  wire  _T_246; 
  wire [31:0] _T_248; 
  wire [32:0] _T_249; 
  wire [32:0] _T_250; 
  wire [32:0] _T_251; 
  wire  _T_252; 
  wire [31:0] _T_253; 
  wire [32:0] _T_254; 
  wire [32:0] _T_255; 
  wire [32:0] _T_256; 
  wire  _T_257; 
  wire  _T_258; 
  wire  _T_261; 
  wire [31:0] _T_264; 
  wire [32:0] _T_265; 
  wire [32:0] _T_266; 
  wire [32:0] _T_267; 
  wire  _T_268; 
  wire  _T_269; 
  wire  _T_273; 
  wire  _T_274; 
  wire  _T_343; 
  wire  _T_360; 
  wire  _T_361; 
  wire  _T_363; 
  wire  _T_364; 
  wire  _T_367; 
  wire  _T_368; 
  wire  _T_370; 
  wire  _T_371; 
  wire  _T_372; 
  wire  _T_374; 
  wire  _T_375; 
  wire [3:0] _T_376; 
  wire  _T_377; 
  wire  _T_379; 
  wire  _T_380; 
  wire  _T_385; 
  wire  _T_515; 
  wire  _T_517; 
  wire  _T_518; 
  wire  _T_528; 
  wire  _T_549; 
  wire  _T_550; 
  wire  _T_553; 
  wire  _T_554; 
  wire  _T_561; 
  wire  _T_563; 
  wire  _T_564; 
  wire  _T_565; 
  wire  _T_567; 
  wire  _T_568; 
  wire  _T_573; 
  wire  _T_588; 
  wire  _T_589; 
  wire  _T_591; 
  wire  _T_599; 
  wire  _T_601; 
  wire  _T_603; 
  wire  _T_604; 
  wire  _T_619; 
  wire [3:0] _T_661; 
  wire [3:0] _T_662; 
  wire  _T_663; 
  wire  _T_665; 
  wire  _T_666; 
  wire  _T_667; 
  wire  _T_669; 
  wire  _T_689; 
  wire  _T_692; 
  wire  _T_693; 
  wire  _T_700; 
  wire  _T_702; 
  wire  _T_703; 
  wire  _T_708; 
  wire  _T_741; 
  wire  _T_743; 
  wire  _T_744; 
  wire  _T_749; 
  wire  _T_795; 
  wire  _T_797; 
  wire  _T_798; 
  wire [2:0] _T_801; 
  wire  _T_802; 
  wire  _T_810; 
  wire  _T_818; 
  wire  _T_826; 
  wire  _T_834; 
  wire  _T_842; 
  wire  _T_850; 
  wire  _T_858; 
  wire  _T_864; 
  wire  _T_865; 
  wire  _T_866; 
  wire  _T_867; 
  wire  _T_868; 
  wire  _T_869; 
  wire  _T_870; 
  wire  _T_871; 
  wire  _T_872; 
  wire  _T_874; 
  wire  _T_875; 
  wire  _T_876; 
  wire  _T_878; 
  wire  _T_879; 
  wire  _T_880; 
  wire  _T_882; 
  wire  _T_883; 
  wire  _T_884; 
  wire  _T_886; 
  wire  _T_887; 
  wire  _T_888; 
  wire  _T_890; 
  wire  _T_891; 
  wire  _T_892; 
  wire  _T_897; 
  wire  _T_898; 
  wire  _T_903; 
  wire  _T_905; 
  wire  _T_906; 
  wire  _T_907; 
  wire  _T_909; 
  wire  _T_910; 
  wire  _T_920; 
  wire  _T_940; 
  wire  _T_942; 
  wire  _T_943; 
  wire  _T_949; 
  wire  _T_966; 
  wire  _T_984; 
  wire [2:0] _T_1521; 
  wire  _T_1522; 
  wire  _T_1530; 
  wire  _T_1538; 
  wire  _T_1546; 
  wire  _T_1554; 
  wire  _T_1562; 
  wire  _T_1570; 
  wire  _T_1578; 
  wire  _T_1584; 
  wire  _T_1585; 
  wire  _T_1586; 
  wire  _T_1587; 
  wire  _T_1588; 
  wire  _T_1589; 
  wire  _T_1590; 
  wire [22:0] _T_1592; 
  wire [7:0] _T_1593; 
  wire [7:0] _T_1594; 
  wire [31:0] _GEN_34; 
  wire [31:0] _T_1595; 
  wire  _T_1596; 
  wire [31:0] _T_1597; 
  wire [32:0] _T_1598; 
  wire [32:0] _T_1599; 
  wire [32:0] _T_1600; 
  wire  _T_1601; 
  wire [31:0] _T_1602; 
  wire [32:0] _T_1603; 
  wire [32:0] _T_1604; 
  wire [32:0] _T_1605; 
  wire  _T_1606; 
  wire [31:0] _T_1607; 
  wire [32:0] _T_1608; 
  wire [32:0] _T_1609; 
  wire [32:0] _T_1610; 
  wire  _T_1611; 
  wire  _T_1613; 
  wire  _T_1614; 
  wire  _T_1745; 
  wire  _T_1747; 
  wire  _T_1748; 
  wire  _T_1750; 
  wire  _T_1751; 
  wire  _T_1752; 
  wire  _T_1754; 
  wire  _T_1755; 
  wire  _T_1757; 
  wire  _T_1758; 
  wire  _T_1759; 
  wire  _T_1761; 
  wire  _T_1762; 
  wire  _T_1767; 
  wire  _T_1785; 
  wire  _T_1800; 
  wire  _T_1808; 
  wire  _T_1812; 
  wire  _T_1813; 
  wire  _T_1882; 
  wire  _T_1899; 
  wire  _T_1900; 
  wire  _T_1911; 
  wire  _T_1913; 
  wire  _T_1914; 
  wire  _T_1919; 
  wire  _T_2049; 
  wire  _T_2059; 
  wire  _T_2061; 
  wire  _T_2062; 
  wire  _T_2067; 
  wire  _T_2081; 
  wire  _T_2099; 
  wire  _T_2101; 
  wire  _T_2102; 
  wire  _T_2103; 
  wire [5:0] _T_2108; 
  wire  _T_2109; 
  wire  _T_2110; 
  reg [5:0] _T_2112; 
  reg [31:0] _RAND_0;
  wire [5:0] _T_2114; 
  wire  _T_2115; 
  reg [2:0] _T_2123; 
  reg [31:0] _RAND_1;
  reg [2:0] _T_2124; 
  reg [31:0] _RAND_2;
  reg [3:0] _T_2125; 
  reg [31:0] _RAND_3;
  reg [5:0] _T_2126; 
  reg [31:0] _RAND_4;
  reg [31:0] _T_2127; 
  reg [31:0] _RAND_5;
  wire  _T_2128; 
  wire  _T_2129; 
  wire  _T_2130; 
  wire  _T_2132; 
  wire  _T_2133; 
  wire  _T_2134; 
  wire  _T_2136; 
  wire  _T_2137; 
  wire  _T_2138; 
  wire  _T_2140; 
  wire  _T_2141; 
  wire  _T_2142; 
  wire  _T_2144; 
  wire  _T_2145; 
  wire  _T_2146; 
  wire  _T_2148; 
  wire  _T_2149; 
  wire  _T_2151; 
  wire  _T_2152; 
  wire [22:0] _T_2154; 
  wire [7:0] _T_2155; 
  wire [7:0] _T_2156; 
  wire [5:0] _T_2157; 
  wire  _T_2158; 
  reg [5:0] _T_2160; 
  reg [31:0] _RAND_6;
  wire [5:0] _T_2162; 
  wire  _T_2163; 
  reg [2:0] _T_2171; 
  reg [31:0] _RAND_7;
  reg [1:0] _T_2172; 
  reg [31:0] _RAND_8;
  reg [3:0] _T_2173; 
  reg [31:0] _RAND_9;
  reg [5:0] _T_2174; 
  reg [31:0] _RAND_10;
  reg  _T_2175; 
  reg [31:0] _RAND_11;
  reg  _T_2176; 
  reg [31:0] _RAND_12;
  wire  _T_2177; 
  wire  _T_2178; 
  wire  _T_2179; 
  wire  _T_2181; 
  wire  _T_2182; 
  wire  _T_2183; 
  wire  _T_2185; 
  wire  _T_2186; 
  wire  _T_2187; 
  wire  _T_2189; 
  wire  _T_2190; 
  wire  _T_2191; 
  wire  _T_2193; 
  wire  _T_2194; 
  wire  _T_2195; 
  wire  _T_2197; 
  wire  _T_2198; 
  wire  _T_2199; 
  wire  _T_2201; 
  wire  _T_2202; 
  wire  _T_2204; 
  wire  _T_2254; 
  wire [5:0] _T_2259; 
  wire  _T_2260; 
  reg [5:0] _T_2262; 
  reg [31:0] _RAND_13;
  wire [5:0] _T_2264; 
  wire  _T_2265; 
  reg [2:0] _T_2273; 
  reg [31:0] _RAND_14;
  reg [2:0] _T_2274; 
  reg [31:0] _RAND_15;
  reg [3:0] _T_2275; 
  reg [31:0] _RAND_16;
  reg [5:0] _T_2276; 
  reg [31:0] _RAND_17;
  reg [31:0] _T_2277; 
  reg [31:0] _RAND_18;
  wire  _T_2278; 
  wire  _T_2279; 
  wire  _T_2280; 
  wire  _T_2282; 
  wire  _T_2283; 
  wire  _T_2284; 
  wire  _T_2286; 
  wire  _T_2287; 
  wire  _T_2288; 
  wire  _T_2290; 
  wire  _T_2291; 
  wire  _T_2292; 
  wire  _T_2294; 
  wire  _T_2295; 
  wire  _T_2296; 
  wire  _T_2298; 
  wire  _T_2299; 
  wire  _T_2301; 
  reg [63:0] _T_2302; 
  reg [63:0] _RAND_19;
  reg [5:0] _T_2312; 
  reg [31:0] _RAND_20;
  wire [5:0] _T_2314; 
  wire  _T_2315; 
  reg [5:0] _T_2331; 
  reg [31:0] _RAND_21;
  wire [5:0] _T_2333; 
  wire  _T_2334; 
  wire  _T_2344; 
  wire [63:0] _T_2346; 
  wire [63:0] _T_2347; 
  wire  _T_2348; 
  wire  _T_2349; 
  wire  _T_2351; 
  wire  _T_2352; 
  wire [63:0] _GEN_27; 
  wire  _T_2356; 
  wire  _T_2358; 
  wire  _T_2359; 
  wire [63:0] _T_2360; 
  wire [63:0] _T_2361; 
  wire [63:0] _T_2362; 
  wire  _T_2363; 
  wire  _T_2365; 
  wire  _T_2366; 
  wire [63:0] _GEN_28; 
  wire  _T_2367; 
  wire  _T_2368; 
  wire  _T_2369; 
  wire  _T_2370; 
  wire  _T_2372; 
  wire  _T_2373; 
  wire [63:0] _T_2374; 
  wire [63:0] _T_2375; 
  wire [63:0] _T_2376; 
  reg [31:0] _T_2377; 
  reg [31:0] _RAND_22;
  wire  _T_2378; 
  wire  _T_2379; 
  wire  _T_2380; 
  wire  _T_2381; 
  wire  _T_2382; 
  wire  _T_2383; 
  wire  _T_2385; 
  wire  _T_2386; 
  wire [31:0] _T_2388; 
  wire  _T_2391; 
  reg  _T_2392; 
  reg [31:0] _RAND_23;
  reg [5:0] _T_2401; 
  reg [31:0] _RAND_24;
  wire [5:0] _T_2403; 
  wire  _T_2404; 
  wire  _T_2414; 
  wire  _T_2415; 
  wire  _T_2416; 
  wire  _T_2417; 
  wire  _T_2418; 
  wire  _T_2419; 
  wire [1:0] _T_2420; 
  wire  _T_2421; 
  wire  _T_2423; 
  wire  _T_2425; 
  wire  _T_2426; 
  wire [1:0] _GEN_31; 
  wire  _T_2428; 
  wire [1:0] _T_2431; 
  wire  _T_2412; 
  wire  _T_2432; 
  wire  _T_2433; 
  wire  _T_2436; 
  wire  _T_2437; 
  wire [1:0] _GEN_32; 
  wire  _T_2438; 
  wire  _T_2427; 
  wire  _T_2439; 
  wire  _T_2440; 
  wire  _GEN_35; 
  wire  _GEN_49; 
  wire  _GEN_65; 
  wire  _GEN_75; 
  wire  _GEN_85; 
  wire  _GEN_95; 
  wire  _GEN_105; 
  wire  _GEN_115; 
  wire  _GEN_123; 
  wire  _GEN_133; 
  wire  _GEN_145; 
  wire  _GEN_157; 
  wire  _GEN_163; 
  wire  _GEN_169; 
  wire  _GEN_175; 
  wire  _GEN_185; 
  wire  _GEN_195; 
  wire  _GEN_207; 
  wire  _GEN_219; 
  wire  _GEN_227; 
  wire  _GEN_235; 
  dual_plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0)) plusarg_reader ( 
    .out(plusarg_reader_out)
  );
  assign _T_7 = io_in_a_bits_source[5:3]; 
  assign _T_8 = _T_7 == 3'h0; 
  assign _T_16 = _T_7 == 3'h1; 
  assign _T_24 = _T_7 == 3'h2; 
  assign _T_32 = _T_7 == 3'h3; 
  assign _T_40 = _T_7 == 3'h4; 
  assign _T_48 = _T_7 == 3'h5; 
  assign _T_56 = _T_7 == 3'h6; 
  assign _T_64 = _T_7 == 3'h7; 
  assign _T_70 = _T_8 | _T_16; 
  assign _T_71 = _T_70 | _T_24; 
  assign _T_72 = _T_71 | _T_32; 
  assign _T_73 = _T_72 | _T_40; 
  assign _T_74 = _T_73 | _T_48; 
  assign _T_75 = _T_74 | _T_56; 
  assign _T_76 = _T_75 | _T_64; 
  assign _T_78 = 23'hff << io_in_a_bits_size; 
  assign _T_79 = _T_78[7:0]; 
  assign _T_80 = ~ _T_79; 
  assign _GEN_33 = {{24'd0}, _T_80}; 
  assign _T_81 = io_in_a_bits_address & _GEN_33; 
  assign _T_82 = _T_81 == 32'h0; 
  assign _T_84 = io_in_a_bits_size[0]; 
  assign _T_85 = 2'h1 << _T_84; 
  assign _T_87 = _T_85 | 2'h1; 
  assign _T_88 = io_in_a_bits_size >= 4'h2; 
  assign _T_89 = _T_87[1]; 
  assign _T_90 = io_in_a_bits_address[1]; 
  assign _T_91 = _T_90 == 1'h0; 
  assign _T_93 = _T_89 & _T_91; 
  assign _T_94 = _T_88 | _T_93; 
  assign _T_96 = _T_89 & _T_90; 
  assign _T_97 = _T_88 | _T_96; 
  assign _T_98 = _T_87[0]; 
  assign _T_99 = io_in_a_bits_address[0]; 
  assign _T_100 = _T_99 == 1'h0; 
  assign _T_101 = _T_91 & _T_100; 
  assign _T_102 = _T_98 & _T_101; 
  assign _T_103 = _T_94 | _T_102; 
  assign _T_104 = _T_91 & _T_99; 
  assign _T_105 = _T_98 & _T_104; 
  assign _T_106 = _T_94 | _T_105; 
  assign _T_107 = _T_90 & _T_100; 
  assign _T_108 = _T_98 & _T_107; 
  assign _T_109 = _T_97 | _T_108; 
  assign _T_110 = _T_90 & _T_99; 
  assign _T_111 = _T_98 & _T_110; 
  assign _T_112 = _T_97 | _T_111; 
  assign _T_115 = {_T_112,_T_109,_T_106,_T_103}; 
  assign _T_246 = io_in_a_bits_opcode == 3'h6; 
  assign _T_248 = io_in_a_bits_address ^ 32'h80000000; 
  assign _T_249 = {1'b0,$signed(_T_248)}; 
  assign _T_250 = $signed(_T_249) & $signed(-33'sh80000000); 
  assign _T_251 = $signed(_T_250); 
  assign _T_252 = $signed(_T_251) == $signed(33'sh0); 
  assign _T_253 = io_in_a_bits_address ^ 32'h40000000; 
  assign _T_254 = {1'b0,$signed(_T_253)}; 
  assign _T_255 = $signed(_T_254) & $signed(-33'sh20000000); 
  assign _T_256 = $signed(_T_255); 
  assign _T_257 = $signed(_T_256) == $signed(33'sh0); 
  assign _T_258 = _T_252 | _T_257; 
  assign _T_261 = io_in_a_bits_size <= 4'h6; 
  assign _T_264 = io_in_a_bits_address ^ 32'h10000000; 
  assign _T_265 = {1'b0,$signed(_T_264)}; 
  assign _T_266 = $signed(_T_265) & $signed(-33'sh10000000); 
  assign _T_267 = $signed(_T_266); 
  assign _T_268 = $signed(_T_267) == $signed(33'sh0); 
  assign _T_269 = _T_261 & _T_268; 
  assign _T_273 = _T_269 | reset; 
  assign _T_274 = _T_273 == 1'h0; 
  assign _T_343 = _T_8 ? _T_261 : 1'h0; 
  assign _T_360 = _T_343 | reset; 
  assign _T_361 = _T_360 == 1'h0; 
  assign _T_363 = _T_76 | reset; 
  assign _T_364 = _T_363 == 1'h0; 
  assign _T_367 = _T_88 | reset; 
  assign _T_368 = _T_367 == 1'h0; 
  assign _T_370 = _T_82 | reset; 
  assign _T_371 = _T_370 == 1'h0; 
  assign _T_372 = io_in_a_bits_param <= 3'h2; 
  assign _T_374 = _T_372 | reset; 
  assign _T_375 = _T_374 == 1'h0; 
  assign _T_376 = ~ io_in_a_bits_mask; 
  assign _T_377 = _T_376 == 4'h0; 
  assign _T_379 = _T_377 | reset; 
  assign _T_380 = _T_379 == 1'h0; 
  assign _T_385 = io_in_a_bits_opcode == 3'h7; 
  assign _T_515 = io_in_a_bits_param != 3'h0; 
  assign _T_517 = _T_515 | reset; 
  assign _T_518 = _T_517 == 1'h0; 
  assign _T_528 = io_in_a_bits_opcode == 3'h4; 
  assign _T_549 = _T_258 | _T_268; 
  assign _T_550 = _T_261 & _T_549; 
  assign _T_553 = _T_550 | reset; 
  assign _T_554 = _T_553 == 1'h0; 
  assign _T_561 = io_in_a_bits_param == 3'h0; 
  assign _T_563 = _T_561 | reset; 
  assign _T_564 = _T_563 == 1'h0; 
  assign _T_565 = io_in_a_bits_mask == _T_115; 
  assign _T_567 = _T_565 | reset; 
  assign _T_568 = _T_567 == 1'h0; 
  assign _T_573 = io_in_a_bits_opcode == 3'h0; 
  assign _T_588 = _T_252 | _T_268; 
  assign _T_589 = _T_261 & _T_588; 
  assign _T_591 = io_in_a_bits_size <= 4'h8; 
  assign _T_599 = _T_591 & _T_257; 
  assign _T_601 = _T_589 | _T_599; 
  assign _T_603 = _T_601 | reset; 
  assign _T_604 = _T_603 == 1'h0; 
  assign _T_619 = io_in_a_bits_opcode == 3'h1; 
  assign _T_661 = ~ _T_115; 
  assign _T_662 = io_in_a_bits_mask & _T_661; 
  assign _T_663 = _T_662 == 4'h0; 
  assign _T_665 = _T_663 | reset; 
  assign _T_666 = _T_665 == 1'h0; 
  assign _T_667 = io_in_a_bits_opcode == 3'h2; 
  assign _T_669 = io_in_a_bits_size <= 4'h3; 
  assign _T_689 = _T_669 & _T_549; 
  assign _T_692 = _T_689 | reset; 
  assign _T_693 = _T_692 == 1'h0; 
  assign _T_700 = io_in_a_bits_param <= 3'h4; 
  assign _T_702 = _T_700 | reset; 
  assign _T_703 = _T_702 == 1'h0; 
  assign _T_708 = io_in_a_bits_opcode == 3'h3; 
  assign _T_741 = io_in_a_bits_param <= 3'h3; 
  assign _T_743 = _T_741 | reset; 
  assign _T_744 = _T_743 == 1'h0; 
  assign _T_749 = io_in_a_bits_opcode == 3'h5; 
  assign _T_795 = io_in_d_bits_opcode <= 3'h6; 
  assign _T_797 = _T_795 | reset; 
  assign _T_798 = _T_797 == 1'h0; 
  assign _T_801 = io_in_d_bits_source[5:3]; 
  assign _T_802 = _T_801 == 3'h0; 
  assign _T_810 = _T_801 == 3'h1; 
  assign _T_818 = _T_801 == 3'h2; 
  assign _T_826 = _T_801 == 3'h3; 
  assign _T_834 = _T_801 == 3'h4; 
  assign _T_842 = _T_801 == 3'h5; 
  assign _T_850 = _T_801 == 3'h6; 
  assign _T_858 = _T_801 == 3'h7; 
  assign _T_864 = _T_802 | _T_810; 
  assign _T_865 = _T_864 | _T_818; 
  assign _T_866 = _T_865 | _T_826; 
  assign _T_867 = _T_866 | _T_834; 
  assign _T_868 = _T_867 | _T_842; 
  assign _T_869 = _T_868 | _T_850; 
  assign _T_870 = _T_869 | _T_858; 
  assign _T_871 = io_in_d_bits_sink < 1'h1; 
  assign _T_872 = io_in_d_bits_opcode == 3'h6; 
  assign _T_874 = _T_870 | reset; 
  assign _T_875 = _T_874 == 1'h0; 
  assign _T_876 = io_in_d_bits_size >= 4'h2; 
  assign _T_878 = _T_876 | reset; 
  assign _T_879 = _T_878 == 1'h0; 
  assign _T_880 = io_in_d_bits_param == 2'h0; 
  assign _T_882 = _T_880 | reset; 
  assign _T_883 = _T_882 == 1'h0; 
  assign _T_884 = io_in_d_bits_corrupt == 1'h0; 
  assign _T_886 = _T_884 | reset; 
  assign _T_887 = _T_886 == 1'h0; 
  assign _T_888 = io_in_d_bits_denied == 1'h0; 
  assign _T_890 = _T_888 | reset; 
  assign _T_891 = _T_890 == 1'h0; 
  assign _T_892 = io_in_d_bits_opcode == 3'h4; 
  assign _T_897 = _T_871 | reset; 
  assign _T_898 = _T_897 == 1'h0; 
  assign _T_903 = io_in_d_bits_param <= 2'h2; 
  assign _T_905 = _T_903 | reset; 
  assign _T_906 = _T_905 == 1'h0; 
  assign _T_907 = io_in_d_bits_param != 2'h2; 
  assign _T_909 = _T_907 | reset; 
  assign _T_910 = _T_909 == 1'h0; 
  assign _T_920 = io_in_d_bits_opcode == 3'h5; 
  assign _T_940 = _T_888 | io_in_d_bits_corrupt; 
  assign _T_942 = _T_940 | reset; 
  assign _T_943 = _T_942 == 1'h0; 
  assign _T_949 = io_in_d_bits_opcode == 3'h0; 
  assign _T_966 = io_in_d_bits_opcode == 3'h1; 
  assign _T_984 = io_in_d_bits_opcode == 3'h2; 
  assign _T_1521 = io_in_c_bits_source[5:3]; 
  assign _T_1522 = _T_1521 == 3'h0; 
  assign _T_1530 = _T_1521 == 3'h1; 
  assign _T_1538 = _T_1521 == 3'h2; 
  assign _T_1546 = _T_1521 == 3'h3; 
  assign _T_1554 = _T_1521 == 3'h4; 
  assign _T_1562 = _T_1521 == 3'h5; 
  assign _T_1570 = _T_1521 == 3'h6; 
  assign _T_1578 = _T_1521 == 3'h7; 
  assign _T_1584 = _T_1522 | _T_1530; 
  assign _T_1585 = _T_1584 | _T_1538; 
  assign _T_1586 = _T_1585 | _T_1546; 
  assign _T_1587 = _T_1586 | _T_1554; 
  assign _T_1588 = _T_1587 | _T_1562; 
  assign _T_1589 = _T_1588 | _T_1570; 
  assign _T_1590 = _T_1589 | _T_1578; 
  assign _T_1592 = 23'hff << io_in_c_bits_size; 
  assign _T_1593 = _T_1592[7:0]; 
  assign _T_1594 = ~ _T_1593; 
  assign _GEN_34 = {{24'd0}, _T_1594}; 
  assign _T_1595 = io_in_c_bits_address & _GEN_34; 
  assign _T_1596 = _T_1595 == 32'h0; 
  assign _T_1597 = io_in_c_bits_address ^ 32'h80000000; 
  assign _T_1598 = {1'b0,$signed(_T_1597)}; 
  assign _T_1599 = $signed(_T_1598) & $signed(-33'sh80000000); 
  assign _T_1600 = $signed(_T_1599); 
  assign _T_1601 = $signed(_T_1600) == $signed(33'sh0); 
  assign _T_1602 = io_in_c_bits_address ^ 32'h40000000; 
  assign _T_1603 = {1'b0,$signed(_T_1602)}; 
  assign _T_1604 = $signed(_T_1603) & $signed(-33'sh20000000); 
  assign _T_1605 = $signed(_T_1604); 
  assign _T_1606 = $signed(_T_1605) == $signed(33'sh0); 
  assign _T_1607 = io_in_c_bits_address ^ 32'h10000000; 
  assign _T_1608 = {1'b0,$signed(_T_1607)}; 
  assign _T_1609 = $signed(_T_1608) & $signed(-33'sh10000000); 
  assign _T_1610 = $signed(_T_1609); 
  assign _T_1611 = $signed(_T_1610) == $signed(33'sh0); 
  assign _T_1613 = _T_1601 | _T_1606; 
  assign _T_1614 = _T_1613 | _T_1611; 
  assign _T_1745 = io_in_c_bits_opcode == 3'h4; 
  assign _T_1747 = _T_1614 | reset; 
  assign _T_1748 = _T_1747 == 1'h0; 
  assign _T_1750 = _T_1590 | reset; 
  assign _T_1751 = _T_1750 == 1'h0; 
  assign _T_1752 = io_in_c_bits_size >= 4'h2; 
  assign _T_1754 = _T_1752 | reset; 
  assign _T_1755 = _T_1754 == 1'h0; 
  assign _T_1757 = _T_1596 | reset; 
  assign _T_1758 = _T_1757 == 1'h0; 
  assign _T_1759 = io_in_c_bits_param <= 3'h5; 
  assign _T_1761 = _T_1759 | reset; 
  assign _T_1762 = _T_1761 == 1'h0; 
  assign _T_1767 = io_in_c_bits_opcode == 3'h5; 
  assign _T_1785 = io_in_c_bits_opcode == 3'h6; 
  assign _T_1800 = io_in_c_bits_size <= 4'h6; 
  assign _T_1808 = _T_1800 & _T_1611; 
  assign _T_1812 = _T_1808 | reset; 
  assign _T_1813 = _T_1812 == 1'h0; 
  assign _T_1882 = _T_1522 ? _T_1800 : 1'h0; 
  assign _T_1899 = _T_1882 | reset; 
  assign _T_1900 = _T_1899 == 1'h0; 
  assign _T_1911 = io_in_c_bits_param <= 3'h2; 
  assign _T_1913 = _T_1911 | reset; 
  assign _T_1914 = _T_1913 == 1'h0; 
  assign _T_1919 = io_in_c_bits_opcode == 3'h7; 
  assign _T_2049 = io_in_c_bits_opcode == 3'h0; 
  assign _T_2059 = io_in_c_bits_param == 3'h0; 
  assign _T_2061 = _T_2059 | reset; 
  assign _T_2062 = _T_2061 == 1'h0; 
  assign _T_2067 = io_in_c_bits_opcode == 3'h1; 
  assign _T_2081 = io_in_c_bits_opcode == 3'h2; 
  assign _T_2099 = io_in_e_bits_sink < 1'h1; 
  assign _T_2101 = _T_2099 | reset; 
  assign _T_2102 = _T_2101 == 1'h0; 
  assign _T_2103 = io_in_a_ready & io_in_a_valid; 
  assign _T_2108 = _T_80[7:2]; 
  assign _T_2109 = io_in_a_bits_opcode[2]; 
  assign _T_2110 = _T_2109 == 1'h0; 
  assign _T_2114 = _T_2112 - 6'h1; 
  assign _T_2115 = _T_2112 == 6'h0; 
  assign _T_2128 = _T_2115 == 1'h0; 
  assign _T_2129 = io_in_a_valid & _T_2128; 
  assign _T_2130 = io_in_a_bits_opcode == _T_2123; 
  assign _T_2132 = _T_2130 | reset; 
  assign _T_2133 = _T_2132 == 1'h0; 
  assign _T_2134 = io_in_a_bits_param == _T_2124; 
  assign _T_2136 = _T_2134 | reset; 
  assign _T_2137 = _T_2136 == 1'h0; 
  assign _T_2138 = io_in_a_bits_size == _T_2125; 
  assign _T_2140 = _T_2138 | reset; 
  assign _T_2141 = _T_2140 == 1'h0; 
  assign _T_2142 = io_in_a_bits_source == _T_2126; 
  assign _T_2144 = _T_2142 | reset; 
  assign _T_2145 = _T_2144 == 1'h0; 
  assign _T_2146 = io_in_a_bits_address == _T_2127; 
  assign _T_2148 = _T_2146 | reset; 
  assign _T_2149 = _T_2148 == 1'h0; 
  assign _T_2151 = _T_2103 & _T_2115; 
  assign _T_2152 = io_in_d_ready & io_in_d_valid; 
  assign _T_2154 = 23'hff << io_in_d_bits_size; 
  assign _T_2155 = _T_2154[7:0]; 
  assign _T_2156 = ~ _T_2155; 
  assign _T_2157 = _T_2156[7:2]; 
  assign _T_2158 = io_in_d_bits_opcode[0]; 
  assign _T_2162 = _T_2160 - 6'h1; 
  assign _T_2163 = _T_2160 == 6'h0; 
  assign _T_2177 = _T_2163 == 1'h0; 
  assign _T_2178 = io_in_d_valid & _T_2177; 
  assign _T_2179 = io_in_d_bits_opcode == _T_2171; 
  assign _T_2181 = _T_2179 | reset; 
  assign _T_2182 = _T_2181 == 1'h0; 
  assign _T_2183 = io_in_d_bits_param == _T_2172; 
  assign _T_2185 = _T_2183 | reset; 
  assign _T_2186 = _T_2185 == 1'h0; 
  assign _T_2187 = io_in_d_bits_size == _T_2173; 
  assign _T_2189 = _T_2187 | reset; 
  assign _T_2190 = _T_2189 == 1'h0; 
  assign _T_2191 = io_in_d_bits_source == _T_2174; 
  assign _T_2193 = _T_2191 | reset; 
  assign _T_2194 = _T_2193 == 1'h0; 
  assign _T_2195 = io_in_d_bits_sink == _T_2175; 
  assign _T_2197 = _T_2195 | reset; 
  assign _T_2198 = _T_2197 == 1'h0; 
  assign _T_2199 = io_in_d_bits_denied == _T_2176; 
  assign _T_2201 = _T_2199 | reset; 
  assign _T_2202 = _T_2201 == 1'h0; 
  assign _T_2204 = _T_2152 & _T_2163; 
  assign _T_2254 = io_in_c_ready & io_in_c_valid; 
  assign _T_2259 = _T_1594[7:2]; 
  assign _T_2260 = io_in_c_bits_opcode[0]; 
  assign _T_2264 = _T_2262 - 6'h1; 
  assign _T_2265 = _T_2262 == 6'h0; 
  assign _T_2278 = _T_2265 == 1'h0; 
  assign _T_2279 = io_in_c_valid & _T_2278; 
  assign _T_2280 = io_in_c_bits_opcode == _T_2273; 
  assign _T_2282 = _T_2280 | reset; 
  assign _T_2283 = _T_2282 == 1'h0; 
  assign _T_2284 = io_in_c_bits_param == _T_2274; 
  assign _T_2286 = _T_2284 | reset; 
  assign _T_2287 = _T_2286 == 1'h0; 
  assign _T_2288 = io_in_c_bits_size == _T_2275; 
  assign _T_2290 = _T_2288 | reset; 
  assign _T_2291 = _T_2290 == 1'h0; 
  assign _T_2292 = io_in_c_bits_source == _T_2276; 
  assign _T_2294 = _T_2292 | reset; 
  assign _T_2295 = _T_2294 == 1'h0; 
  assign _T_2296 = io_in_c_bits_address == _T_2277; 
  assign _T_2298 = _T_2296 | reset; 
  assign _T_2299 = _T_2298 == 1'h0; 
  assign _T_2301 = _T_2254 & _T_2265; 
  assign _T_2314 = _T_2312 - 6'h1; 
  assign _T_2315 = _T_2312 == 6'h0; 
  assign _T_2333 = _T_2331 - 6'h1; 
  assign _T_2334 = _T_2331 == 6'h0; 
  assign _T_2344 = _T_2103 & _T_2315; 
  assign _T_2346 = 64'h1 << io_in_a_bits_source; 
  assign _T_2347 = _T_2302 >> io_in_a_bits_source; 
  assign _T_2348 = _T_2347[0]; 
  assign _T_2349 = _T_2348 == 1'h0; 
  assign _T_2351 = _T_2349 | reset; 
  assign _T_2352 = _T_2351 == 1'h0; 
  assign _GEN_27 = _T_2344 ? _T_2346 : 64'h0; 
  assign _T_2356 = _T_2152 & _T_2334; 
  assign _T_2358 = _T_872 == 1'h0; 
  assign _T_2359 = _T_2356 & _T_2358; 
  assign _T_2360 = 64'h1 << io_in_d_bits_source; 
  assign _T_2361 = _GEN_27 | _T_2302; 
  assign _T_2362 = _T_2361 >> io_in_d_bits_source; 
  assign _T_2363 = _T_2362[0]; 
  assign _T_2365 = _T_2363 | reset; 
  assign _T_2366 = _T_2365 == 1'h0; 
  assign _GEN_28 = _T_2359 ? _T_2360 : 64'h0; 
  assign _T_2367 = _GEN_27 != _GEN_28; 
  assign _T_2368 = _GEN_27 != 64'h0; 
  assign _T_2369 = _T_2368 == 1'h0; 
  assign _T_2370 = _T_2367 | _T_2369; 
  assign _T_2372 = _T_2370 | reset; 
  assign _T_2373 = _T_2372 == 1'h0; 
  assign _T_2374 = _T_2302 | _GEN_27; 
  assign _T_2375 = ~ _GEN_28; 
  assign _T_2376 = _T_2374 & _T_2375; 
  assign _T_2378 = _T_2302 != 64'h0; 
  assign _T_2379 = _T_2378 == 1'h0; 
  assign _T_2380 = plusarg_reader_out == 32'h0; 
  assign _T_2381 = _T_2379 | _T_2380; 
  assign _T_2382 = _T_2377 < plusarg_reader_out; 
  assign _T_2383 = _T_2381 | _T_2382; 
  assign _T_2385 = _T_2383 | reset; 
  assign _T_2386 = _T_2385 == 1'h0; 
  assign _T_2388 = _T_2377 + 32'h1; 
  assign _T_2391 = _T_2103 | _T_2152; 
  assign _T_2403 = _T_2401 - 6'h1; 
  assign _T_2404 = _T_2401 == 6'h0; 
  assign _T_2414 = _T_2152 & _T_2404; 
  assign _T_2415 = io_in_d_bits_opcode[2]; 
  assign _T_2416 = io_in_d_bits_opcode[1]; 
  assign _T_2417 = _T_2416 == 1'h0; 
  assign _T_2418 = _T_2415 & _T_2417; 
  assign _T_2419 = _T_2414 & _T_2418; 
  assign _T_2420 = 2'h1 << io_in_d_bits_sink; 
  assign _T_2421 = _T_2392 >> io_in_d_bits_sink; 
  assign _T_2423 = _T_2421 == 1'h0; 
  assign _T_2425 = _T_2423 | reset; 
  assign _T_2426 = _T_2425 == 1'h0; 
  assign _GEN_31 = _T_2419 ? _T_2420 : 2'h0; 
  assign _T_2428 = io_in_e_ready & io_in_e_valid; 
  assign _T_2431 = 2'h1 << io_in_e_bits_sink; 
  assign _T_2412 = _GEN_31[0]; 
  assign _T_2432 = _T_2412 | _T_2392; 
  assign _T_2433 = _T_2432 >> io_in_e_bits_sink; 
  assign _T_2436 = _T_2433 | reset; 
  assign _T_2437 = _T_2436 == 1'h0; 
  assign _GEN_32 = _T_2428 ? _T_2431 : 2'h0; 
  assign _T_2438 = _T_2392 | _T_2412; 
  assign _T_2427 = _GEN_32[0]; 
  assign _T_2439 = ~ _T_2427; 
  assign _T_2440 = _T_2438 & _T_2439; 
  assign _GEN_35 = io_in_a_valid & _T_246; 
  assign _GEN_49 = io_in_a_valid & _T_385; 
  assign _GEN_65 = io_in_a_valid & _T_528; 
  assign _GEN_75 = io_in_a_valid & _T_573; 
  assign _GEN_85 = io_in_a_valid & _T_619; 
  assign _GEN_95 = io_in_a_valid & _T_667; 
  assign _GEN_105 = io_in_a_valid & _T_708; 
  assign _GEN_115 = io_in_a_valid & _T_749; 
  assign _GEN_123 = io_in_d_valid & _T_872; 
  assign _GEN_133 = io_in_d_valid & _T_892; 
  assign _GEN_145 = io_in_d_valid & _T_920; 
  assign _GEN_157 = io_in_d_valid & _T_949; 
  assign _GEN_163 = io_in_d_valid & _T_966; 
  assign _GEN_169 = io_in_d_valid & _T_984; 
  assign _GEN_175 = io_in_c_valid & _T_1745; 
  assign _GEN_185 = io_in_c_valid & _T_1767; 
  assign _GEN_195 = io_in_c_valid & _T_1785; 
  assign _GEN_207 = io_in_c_valid & _T_1919; 
  assign _GEN_219 = io_in_c_valid & _T_2049; 
  assign _GEN_227 = io_in_c_valid & _T_2067; 
  assign _GEN_235 = io_in_c_valid & _T_2081; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2112 = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_2123 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2124 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_2125 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_2126 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_2127 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_2160 = _RAND_6[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_2171 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_2172 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_2173 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_2174 = _RAND_10[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_2175 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_2176 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_2262 = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_2273 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_2274 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_2275 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_2276 = _RAND_17[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_2277 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  _T_2302 = _RAND_19[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_2312 = _RAND_20[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_2331 = _RAND_21[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_2377 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_2392 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_2401 = _RAND_24[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_2112 <= 6'h0;
    end else begin
      if (_T_2103) begin
        if (_T_2115) begin
          if (_T_2110) begin
            _T_2112 <= _T_2108;
          end else begin
            _T_2112 <= 6'h0;
          end
        end else begin
          _T_2112 <= _T_2114;
        end
      end
    end
    if (_T_2151) begin
      _T_2123 <= io_in_a_bits_opcode;
    end
    if (_T_2151) begin
      _T_2124 <= io_in_a_bits_param;
    end
    if (_T_2151) begin
      _T_2125 <= io_in_a_bits_size;
    end
    if (_T_2151) begin
      _T_2126 <= io_in_a_bits_source;
    end
    if (_T_2151) begin
      _T_2127 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_2160 <= 6'h0;
    end else begin
      if (_T_2152) begin
        if (_T_2163) begin
          if (_T_2158) begin
            _T_2160 <= _T_2157;
          end else begin
            _T_2160 <= 6'h0;
          end
        end else begin
          _T_2160 <= _T_2162;
        end
      end
    end
    if (_T_2204) begin
      _T_2171 <= io_in_d_bits_opcode;
    end
    if (_T_2204) begin
      _T_2172 <= io_in_d_bits_param;
    end
    if (_T_2204) begin
      _T_2173 <= io_in_d_bits_size;
    end
    if (_T_2204) begin
      _T_2174 <= io_in_d_bits_source;
    end
    if (_T_2204) begin
      _T_2175 <= io_in_d_bits_sink;
    end
    if (_T_2204) begin
      _T_2176 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_2262 <= 6'h0;
    end else begin
      if (_T_2254) begin
        if (_T_2265) begin
          if (_T_2260) begin
            _T_2262 <= _T_2259;
          end else begin
            _T_2262 <= 6'h0;
          end
        end else begin
          _T_2262 <= _T_2264;
        end
      end
    end
    if (_T_2301) begin
      _T_2273 <= io_in_c_bits_opcode;
    end
    if (_T_2301) begin
      _T_2274 <= io_in_c_bits_param;
    end
    if (_T_2301) begin
      _T_2275 <= io_in_c_bits_size;
    end
    if (_T_2301) begin
      _T_2276 <= io_in_c_bits_source;
    end
    if (_T_2301) begin
      _T_2277 <= io_in_c_bits_address;
    end
    if (reset) begin
      _T_2302 <= 64'h0;
    end else begin
      _T_2302 <= _T_2376;
    end
    if (reset) begin
      _T_2312 <= 6'h0;
    end else begin
      if (_T_2103) begin
        if (_T_2315) begin
          if (_T_2110) begin
            _T_2312 <= _T_2108;
          end else begin
            _T_2312 <= 6'h0;
          end
        end else begin
          _T_2312 <= _T_2314;
        end
      end
    end
    if (reset) begin
      _T_2331 <= 6'h0;
    end else begin
      if (_T_2152) begin
        if (_T_2334) begin
          if (_T_2158) begin
            _T_2331 <= _T_2157;
          end else begin
            _T_2331 <= 6'h0;
          end
        end else begin
          _T_2331 <= _T_2333;
        end
      end
    end
    if (reset) begin
      _T_2377 <= 32'h0;
    end else begin
      if (_T_2391) begin
        _T_2377 <= 32'h0;
      end else begin
        _T_2377 <= _T_2388;
      end
    end
    if (reset) begin
      _T_2392 <= 1'h0;
    end else begin
      _T_2392 <= _T_2440;
    end
    if (reset) begin
      _T_2401 <= 6'h0;
    end else begin
      if (_T_2152) begin
        if (_T_2404) begin
          if (_T_2158) begin
            _T_2401 <= _T_2157;
          end else begin
            _T_2401 <= 6'h0;
          end
        end else begin
          _T_2401 <= _T_2403;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel has invalid opcode (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:39 assert (TLMessages.isA(bundle.opcode), \"'A' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:46 assert (visible(edge.address(bundle), bundle.source, edge), \"'A' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_274) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_274) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_361) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_361) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_364) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_364) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_368) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_368) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_371) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_371) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_375) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_375) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_380) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_380) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:56 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_274) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_274) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_361) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_361) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_364) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_364) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_368) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_368) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_371) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_371) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_375) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_375) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_518) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_518) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_380) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_380) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:68 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_554) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_554) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_364) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_364) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_371) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_371) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_564) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_564) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_568) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_568) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:77 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_604) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_604) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_364) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_364) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_371) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_371) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_564) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_564) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_568) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_568) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_604) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_604) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_364) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_364) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_371) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_371) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_564) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_564) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_666) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_666) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_693) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_693) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_364) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_364) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_371) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_371) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_703) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_703) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_568) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_568) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_693) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_693) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_364) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_364) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_371) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_371) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_744) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_744) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_568) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_568) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_604) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_604) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_364) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_364) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_371) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_371) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_568) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_568) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:117 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_798) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_798) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_875) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_875) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_879) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_879) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_883) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_883) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_887) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_887) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_891) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_891) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_875) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_875) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_898) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:285 assert (sink_ok, \"'D' channel Grant carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_898) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_879) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_879) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_906) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_906) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_910) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_910) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_887) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_887) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is denied (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:290 assert (deny_put_ok || !bundle.denied, \"'D' channel Grant is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_875) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_875) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_898) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:295 assert (sink_ok, \"'D' channel GrantData carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_898) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_879) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_879) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_906) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_906) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_910) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_910) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_145 & _T_943) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_145 & _T_943) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:300 assert (deny_get_ok || !bundle.denied, \"'D' channel GrantData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_157 & _T_875) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_157 & _T_875) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_157 & _T_883) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_157 & _T_883) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_157 & _T_887) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_157 & _T_887) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is denied (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:308 assert (deny_put_ok || !bundle.denied, \"'D' channel AccessAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_875) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_875) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_883) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_883) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_943) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_943) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:316 assert (deny_get_ok || !bundle.denied, \"'D' channel AccessAckData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_169 & _T_875) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_169 & _T_875) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_169 & _T_883) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_169 & _T_883) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_169 & _T_887) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_169 & _T_887) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is denied (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:324 assert (deny_put_ok || !bundle.denied, \"'D' channel HintAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel has invalid opcode (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:122 assert (TLMessages.isB(bundle.opcode), \"'B' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:124 assert (visible(edge.address(bundle), bundle.source, edge), \"'B' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Probe type unsupported by client (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:133 assert (edge.client.supportsProbe(bundle.source, bundle.size), \"'B' channel carries Probe type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:134 assert (address_ok, \"'B' channel Probe carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries source that is not first source (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:135 assert (legal_source, \"'B' channel Probe carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:136 assert (is_aligned, \"'B' channel Probe address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:137 assert (TLPermissions.isCap(bundle.param), \"'B' channel Probe carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe contains invalid mask (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:138 assert (bundle.mask === mask, \"'B' channel Probe contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe is corrupt (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:139 assert (!bundle.corrupt, \"'B' channel Probe is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Get type unsupported by client (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:143 assert (edge.client.supportsGet(bundle.source, bundle.size), \"'B' channel carries Get type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries unmanaged address (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:144 assert (address_ok, \"'B' channel Get carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries source that is not first source (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:145 assert (legal_source, \"'B' channel Get carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:146 assert (is_aligned, \"'B' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries invalid param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:147 assert (bundle.param === UInt(0), \"'B' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get contains invalid mask (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:148 assert (bundle.mask === mask, \"'B' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get is corrupt (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:149 assert (!bundle.corrupt, \"'B' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutFull type unsupported by client (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:153 assert (edge.client.supportsPutFull(bundle.source, bundle.size), \"'B' channel carries PutFull type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries unmanaged address (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:154 assert (address_ok, \"'B' channel PutFull carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries source that is not first source (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:155 assert (legal_source, \"'B' channel PutFull carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:156 assert (is_aligned, \"'B' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries invalid param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:157 assert (bundle.param === UInt(0), \"'B' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull contains invalid mask (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:158 assert (bundle.mask === mask, \"'B' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutPartial type unsupported by client (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:162 assert (edge.client.supportsPutPartial(bundle.source, bundle.size), \"'B' channel carries PutPartial type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:163 assert (address_ok, \"'B' channel PutPartial carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:164 assert (legal_source, \"'B' channel PutPartial carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:165 assert (is_aligned, \"'B' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries invalid param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:166 assert (bundle.param === UInt(0), \"'B' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial contains invalid mask (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:167 assert ((bundle.mask & ~mask) === UInt(0), \"'B' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Arithmetic type unsupported by client (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:171 assert (edge.client.supportsArithmetic(bundle.source, bundle.size), \"'B' channel carries Arithmetic type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:172 assert (address_ok, \"'B' channel Arithmetic carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:173 assert (legal_source, \"'B' channel Arithmetic carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:174 assert (is_aligned, \"'B' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries invalid opcode param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:175 assert (TLAtomics.isArithmetic(bundle.param), \"'B' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:176 assert (bundle.mask === mask, \"'B' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Logical type unsupported by client (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:180 assert (edge.client.supportsLogical(bundle.source, bundle.size), \"'B' channel carries Logical type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries unmanaged address (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:181 assert (address_ok, \"'B' channel Logical carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries source that is not first source (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:182 assert (legal_source, \"'B' channel Logical carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:183 assert (is_aligned, \"'B' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries invalid opcode param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:184 assert (TLAtomics.isLogical(bundle.param), \"'B' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical contains invalid mask (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:185 assert (bundle.mask === mask, \"'B' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Hint type unsupported by client (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:189 assert (edge.client.supportsHint(bundle.source, bundle.size), \"'B' channel carries Hint type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries unmanaged address (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:190 assert (address_ok, \"'B' channel Hint carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries source that is not first source (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:191 assert (legal_source, \"'B' channel Hint carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:192 assert (is_aligned, \"'B' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint contains invalid mask (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:193 assert (bundle.mask === mask, \"'B' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint is corrupt (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:194 assert (!bundle.corrupt, \"'B' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel has invalid opcode (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:199 assert (TLMessages.isC(bundle.opcode), \"'C' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:205 assert (visible(edge.address(bundle), bundle.source, edge), \"'C' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1748) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:208 assert (address_ok, \"'C' channel ProbeAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1748) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1751) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:209 assert (source_ok, \"'C' channel ProbeAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1751) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1755) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:210 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1755) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1758) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:211 assert (is_aligned, \"'C' channel ProbeAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1758) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_1762) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:212 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAck carries invalid report param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_175 & _T_1762) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck is corrupt (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:213 assert (!bundle.corrupt, \"'C' channel ProbeAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & _T_1748) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:217 assert (address_ok, \"'C' channel ProbeAckData carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & _T_1748) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & _T_1751) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:218 assert (source_ok, \"'C' channel ProbeAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & _T_1751) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & _T_1755) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:219 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAckData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & _T_1755) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & _T_1758) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:220 assert (is_aligned, \"'C' channel ProbeAckData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & _T_1758) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & _T_1762) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:221 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAckData carries invalid report param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & _T_1762) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1813) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:225 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries Release type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1813) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1900) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:226 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1900) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1751) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:227 assert (source_ok, \"'C' channel Release carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1751) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1755) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:228 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel Release smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1755) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1758) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:229 assert (is_aligned, \"'C' channel Release address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1758) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1914) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid shrink param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:230 assert (TLPermissions.isShrink(bundle.param), \"'C' channel Release carries invalid shrink param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1914) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release is corrupt (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:231 assert (!bundle.corrupt, \"'C' channel Release is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_207 & _T_1813) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:235 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries ReleaseData type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_207 & _T_1813) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_207 & _T_1900) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:236 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_207 & _T_1900) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_207 & _T_1751) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:237 assert (source_ok, \"'C' channel ReleaseData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_207 & _T_1751) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_207 & _T_1755) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:238 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ReleaseData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_207 & _T_1755) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_207 & _T_1758) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:239 assert (is_aligned, \"'C' channel ReleaseData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_207 & _T_1758) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_207 & _T_1914) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid shrink param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:240 assert (TLPermissions.isShrink(bundle.param), \"'C' channel ReleaseData carries invalid shrink param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_207 & _T_1914) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1748) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:244 assert (address_ok, \"'C' channel AccessAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1748) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1751) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:245 assert (source_ok, \"'C' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1751) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1758) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:246 assert (is_aligned, \"'C' channel AccessAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1758) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_2062) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:247 assert (bundle.param === UInt(0), \"'C' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_2062) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck is corrupt (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:248 assert (!bundle.corrupt, \"'C' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_227 & _T_1748) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:252 assert (address_ok, \"'C' channel AccessAckData carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_227 & _T_1748) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_227 & _T_1751) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:253 assert (source_ok, \"'C' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_227 & _T_1751) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_227 & _T_1758) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:254 assert (is_aligned, \"'C' channel AccessAckData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_227 & _T_1758) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_227 & _T_2062) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:255 assert (bundle.param === UInt(0), \"'C' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_227 & _T_2062) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_235 & _T_1748) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:259 assert (address_ok, \"'C' channel HintAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_1748) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_235 & _T_1751) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:260 assert (source_ok, \"'C' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_1751) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_235 & _T_1758) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:261 assert (is_aligned, \"'C' channel HintAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_1758) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_235 & _T_2062) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:262 assert (bundle.param === UInt(0), \"'C' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_2062) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck is corrupt (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:263 assert (!bundle.corrupt, \"'C' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_e_valid & _T_2102) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channels carries invalid sink ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:330 assert (sink_ok, \"'E' channels carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_e_valid & _T_2102) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2129 & _T_2133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2129 & _T_2133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2129 & _T_2137) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2129 & _T_2137) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2129 & _T_2141) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2129 & _T_2141) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2129 & _T_2145) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2129 & _T_2145) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2129 & _T_2149) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2129 & _T_2149) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2178 & _T_2182) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2178 & _T_2182) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2178 & _T_2186) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2178 & _T_2186) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2178 & _T_2190) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2178 & _T_2190) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2178 & _T_2194) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2178 & _T_2194) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2178 & _T_2198) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2178 & _T_2198) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2178 & _T_2202) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2178 & _T_2202) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel opcode changed within multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:378 assert (b.bits.opcode === opcode, \"'B' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:379 assert (b.bits.param  === param,  \"'B' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel size changed within multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:380 assert (b.bits.size   === size,   \"'B' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel source changed within multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:381 assert (b.bits.source === source, \"'B' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:382 assert (b.bits.address=== address,\"'B' channel addresss changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2279 & _T_2283) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:401 assert (c.bits.opcode === opcode, \"'C' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2279 & _T_2283) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2279 & _T_2287) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:402 assert (c.bits.param  === param,  \"'C' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2279 & _T_2287) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2279 & _T_2291) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:403 assert (c.bits.size   === size,   \"'C' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2279 & _T_2291) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2279 & _T_2295) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:404 assert (c.bits.source === source, \"'C' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2279 & _T_2295) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2279 & _T_2299) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:405 assert (c.bits.address=== address,\"'C' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2279 & _T_2299) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2344 & _T_2352) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2344 & _T_2352) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2359 & _T_2366) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2359 & _T_2366) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2373) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2373) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2386) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:479 assert (!inflight.orR || limit === UInt(0) || watchdog < limit, \"TileLink timeout expired\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2386) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2419 & _T_2426) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:494 assert(!inflight(bundle.d.bits.sink), \"'D' channel re-used a sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2419 & _T_2426) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2428 & _T_2437) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at dual_ChipLink.scala:78:16)\n    at Monitor.scala:500 assert((d_set | inflight)(bundle.e.bits.sink), \"'E' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2428 & _T_2437) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLMonitor_7( 
  input        clock, 
  input        reset, 
  input        io_in_d_valid, 
  input  [2:0] io_in_d_bits_opcode, 
  input  [1:0] io_in_d_bits_param, 
  input  [3:0] io_in_d_bits_size, 
  input        io_in_d_bits_source, 
  input        io_in_d_bits_sink, 
  input        io_in_d_bits_denied, 
  input        io_in_d_bits_corrupt 
);
  wire [31:0] plusarg_reader_out; 
  wire  _T_444; 
  wire  _T_446; 
  wire  _T_447; 
  wire  _T_448; 
  wire  _T_450; 
  wire  _T_451; 
  wire  _T_453; 
  wire  _T_454; 
  wire  _T_455; 
  wire  _T_457; 
  wire  _T_458; 
  wire  _T_459; 
  wire  _T_461; 
  wire  _T_462; 
  wire  _T_463; 
  wire  _T_465; 
  wire  _T_466; 
  wire  _T_467; 
  wire  _T_469; 
  wire  _T_470; 
  wire  _T_471; 
  wire  _T_476; 
  wire  _T_477; 
  wire  _T_482; 
  wire  _T_484; 
  wire  _T_485; 
  wire  _T_486; 
  wire  _T_488; 
  wire  _T_489; 
  wire  _T_499; 
  wire  _T_519; 
  wire  _T_521; 
  wire  _T_522; 
  wire  _T_528; 
  wire  _T_545; 
  wire  _T_563; 
  wire [22:0] _T_1103; 
  wire [7:0] _T_1104; 
  wire [7:0] _T_1105; 
  wire [5:0] _T_1106; 
  wire  _T_1107; 
  reg [5:0] _T_1109; 
  reg [31:0] _RAND_0;
  wire [5:0] _T_1111; 
  wire  _T_1112; 
  reg [2:0] _T_1120; 
  reg [31:0] _RAND_1;
  reg [1:0] _T_1121; 
  reg [31:0] _RAND_2;
  reg [3:0] _T_1122; 
  reg [31:0] _RAND_3;
  reg  _T_1123; 
  reg [31:0] _RAND_4;
  reg  _T_1124; 
  reg [31:0] _RAND_5;
  reg  _T_1125; 
  reg [31:0] _RAND_6;
  wire  _T_1126; 
  wire  _T_1127; 
  wire  _T_1128; 
  wire  _T_1130; 
  wire  _T_1131; 
  wire  _T_1132; 
  wire  _T_1134; 
  wire  _T_1135; 
  wire  _T_1136; 
  wire  _T_1138; 
  wire  _T_1139; 
  wire  _T_1140; 
  wire  _T_1142; 
  wire  _T_1143; 
  wire  _T_1144; 
  wire  _T_1146; 
  wire  _T_1147; 
  wire  _T_1148; 
  wire  _T_1150; 
  wire  _T_1151; 
  wire  _T_1153; 
  reg  _T_1251; 
  reg [31:0] _RAND_7;
  reg [5:0] _T_1280; 
  reg [31:0] _RAND_8;
  wire [5:0] _T_1282; 
  wire  _T_1283; 
  wire  _T_1298; 
  wire  _T_1305; 
  wire  _T_1307; 
  wire  _T_1308; 
  wire [1:0] _T_1309; 
  wire  _T_1311; 
  wire  _T_1314; 
  wire  _T_1315; 
  wire [1:0] _GEN_28; 
  wire  _T_1302; 
  wire  _T_1324; 
  wire  _T_1325; 
  reg [31:0] _T_1326; 
  reg [31:0] _RAND_9;
  wire  _T_1329; 
  wire  _T_1330; 
  wire  _T_1331; 
  wire  _T_1332; 
  wire  _T_1334; 
  wire  _T_1335; 
  wire [31:0] _T_1337; 
  reg  _T_1341; 
  reg [31:0] _RAND_10;
  reg [5:0] _T_1350; 
  reg [31:0] _RAND_11;
  wire [5:0] _T_1352; 
  wire  _T_1353; 
  wire  _T_1363; 
  wire  _T_1364; 
  wire  _T_1365; 
  wire  _T_1366; 
  wire  _T_1367; 
  wire  _T_1368; 
  wire [1:0] _T_1369; 
  wire  _T_1370; 
  wire  _T_1372; 
  wire  _T_1374; 
  wire  _T_1375; 
  wire [1:0] _GEN_31; 
  wire  _T_1361; 
  wire  _T_1387; 
  wire  _GEN_33; 
  wire  _GEN_43; 
  wire  _GEN_55; 
  wire  _GEN_67; 
  wire  _GEN_73; 
  wire  _GEN_79; 
  dual_plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0)) plusarg_reader ( 
    .out(plusarg_reader_out)
  );
  assign _T_444 = io_in_d_bits_opcode <= 3'h6; 
  assign _T_446 = _T_444 | reset; 
  assign _T_447 = _T_446 == 1'h0; 
  assign _T_448 = io_in_d_bits_source == 1'h0; 
  assign _T_450 = io_in_d_bits_sink < 1'h1; 
  assign _T_451 = io_in_d_bits_opcode == 3'h6; 
  assign _T_453 = _T_448 | reset; 
  assign _T_454 = _T_453 == 1'h0; 
  assign _T_455 = io_in_d_bits_size >= 4'h2; 
  assign _T_457 = _T_455 | reset; 
  assign _T_458 = _T_457 == 1'h0; 
  assign _T_459 = io_in_d_bits_param == 2'h0; 
  assign _T_461 = _T_459 | reset; 
  assign _T_462 = _T_461 == 1'h0; 
  assign _T_463 = io_in_d_bits_corrupt == 1'h0; 
  assign _T_465 = _T_463 | reset; 
  assign _T_466 = _T_465 == 1'h0; 
  assign _T_467 = io_in_d_bits_denied == 1'h0; 
  assign _T_469 = _T_467 | reset; 
  assign _T_470 = _T_469 == 1'h0; 
  assign _T_471 = io_in_d_bits_opcode == 3'h4; 
  assign _T_476 = _T_450 | reset; 
  assign _T_477 = _T_476 == 1'h0; 
  assign _T_482 = io_in_d_bits_param <= 2'h2; 
  assign _T_484 = _T_482 | reset; 
  assign _T_485 = _T_484 == 1'h0; 
  assign _T_486 = io_in_d_bits_param != 2'h2; 
  assign _T_488 = _T_486 | reset; 
  assign _T_489 = _T_488 == 1'h0; 
  assign _T_499 = io_in_d_bits_opcode == 3'h5; 
  assign _T_519 = _T_467 | io_in_d_bits_corrupt; 
  assign _T_521 = _T_519 | reset; 
  assign _T_522 = _T_521 == 1'h0; 
  assign _T_528 = io_in_d_bits_opcode == 3'h0; 
  assign _T_545 = io_in_d_bits_opcode == 3'h1; 
  assign _T_563 = io_in_d_bits_opcode == 3'h2; 
  assign _T_1103 = 23'hff << io_in_d_bits_size; 
  assign _T_1104 = _T_1103[7:0]; 
  assign _T_1105 = ~ _T_1104; 
  assign _T_1106 = _T_1105[7:2]; 
  assign _T_1107 = io_in_d_bits_opcode[0]; 
  assign _T_1111 = _T_1109 - 6'h1; 
  assign _T_1112 = _T_1109 == 6'h0; 
  assign _T_1126 = _T_1112 == 1'h0; 
  assign _T_1127 = io_in_d_valid & _T_1126; 
  assign _T_1128 = io_in_d_bits_opcode == _T_1120; 
  assign _T_1130 = _T_1128 | reset; 
  assign _T_1131 = _T_1130 == 1'h0; 
  assign _T_1132 = io_in_d_bits_param == _T_1121; 
  assign _T_1134 = _T_1132 | reset; 
  assign _T_1135 = _T_1134 == 1'h0; 
  assign _T_1136 = io_in_d_bits_size == _T_1122; 
  assign _T_1138 = _T_1136 | reset; 
  assign _T_1139 = _T_1138 == 1'h0; 
  assign _T_1140 = io_in_d_bits_source == _T_1123; 
  assign _T_1142 = _T_1140 | reset; 
  assign _T_1143 = _T_1142 == 1'h0; 
  assign _T_1144 = io_in_d_bits_sink == _T_1124; 
  assign _T_1146 = _T_1144 | reset; 
  assign _T_1147 = _T_1146 == 1'h0; 
  assign _T_1148 = io_in_d_bits_denied == _T_1125; 
  assign _T_1150 = _T_1148 | reset; 
  assign _T_1151 = _T_1150 == 1'h0; 
  assign _T_1153 = io_in_d_valid & _T_1112; 
  assign _T_1282 = _T_1280 - 6'h1; 
  assign _T_1283 = _T_1280 == 6'h0; 
  assign _T_1298 = _T_1251 == 1'h0; 
  assign _T_1305 = io_in_d_valid & _T_1283; 
  assign _T_1307 = _T_451 == 1'h0; 
  assign _T_1308 = _T_1305 & _T_1307; 
  assign _T_1309 = 2'h1 << io_in_d_bits_source; 
  assign _T_1311 = _T_1251 >> io_in_d_bits_source; 
  assign _T_1314 = _T_1311 | reset; 
  assign _T_1315 = _T_1314 == 1'h0; 
  assign _GEN_28 = _T_1308 ? _T_1309 : 2'h0; 
  assign _T_1302 = _GEN_28[0]; 
  assign _T_1324 = ~ _T_1302; 
  assign _T_1325 = _T_1251 & _T_1324; 
  assign _T_1329 = plusarg_reader_out == 32'h0; 
  assign _T_1330 = _T_1298 | _T_1329; 
  assign _T_1331 = _T_1326 < plusarg_reader_out; 
  assign _T_1332 = _T_1330 | _T_1331; 
  assign _T_1334 = _T_1332 | reset; 
  assign _T_1335 = _T_1334 == 1'h0; 
  assign _T_1337 = _T_1326 + 32'h1; 
  assign _T_1352 = _T_1350 - 6'h1; 
  assign _T_1353 = _T_1350 == 6'h0; 
  assign _T_1363 = io_in_d_valid & _T_1353; 
  assign _T_1364 = io_in_d_bits_opcode[2]; 
  assign _T_1365 = io_in_d_bits_opcode[1]; 
  assign _T_1366 = _T_1365 == 1'h0; 
  assign _T_1367 = _T_1364 & _T_1366; 
  assign _T_1368 = _T_1363 & _T_1367; 
  assign _T_1369 = 2'h1 << io_in_d_bits_sink; 
  assign _T_1370 = _T_1341 >> io_in_d_bits_sink; 
  assign _T_1372 = _T_1370 == 1'h0; 
  assign _T_1374 = _T_1372 | reset; 
  assign _T_1375 = _T_1374 == 1'h0; 
  assign _GEN_31 = _T_1368 ? _T_1369 : 2'h0; 
  assign _T_1361 = _GEN_31[0]; 
  assign _T_1387 = _T_1341 | _T_1361; 
  assign _GEN_33 = io_in_d_valid & _T_451; 
  assign _GEN_43 = io_in_d_valid & _T_471; 
  assign _GEN_55 = io_in_d_valid & _T_499; 
  assign _GEN_67 = io_in_d_valid & _T_528; 
  assign _GEN_73 = io_in_d_valid & _T_545; 
  assign _GEN_79 = io_in_d_valid & _T_563; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1109 = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1120 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1121 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1122 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1123 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1124 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_1125 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_1251 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1280 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_1326 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_1341 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_1350 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_1109 <= 6'h0;
    end else begin
      if (io_in_d_valid) begin
        if (_T_1112) begin
          if (_T_1107) begin
            _T_1109 <= _T_1106;
          end else begin
            _T_1109 <= 6'h0;
          end
        end else begin
          _T_1109 <= _T_1111;
        end
      end
    end
    if (_T_1153) begin
      _T_1120 <= io_in_d_bits_opcode;
    end
    if (_T_1153) begin
      _T_1121 <= io_in_d_bits_param;
    end
    if (_T_1153) begin
      _T_1122 <= io_in_d_bits_size;
    end
    if (_T_1153) begin
      _T_1123 <= io_in_d_bits_source;
    end
    if (_T_1153) begin
      _T_1124 <= io_in_d_bits_sink;
    end
    if (_T_1153) begin
      _T_1125 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_1251 <= 1'h0;
    end else begin
      _T_1251 <= _T_1325;
    end
    if (reset) begin
      _T_1280 <= 6'h0;
    end else begin
      if (io_in_d_valid) begin
        if (_T_1283) begin
          if (_T_1107) begin
            _T_1280 <= _T_1106;
          end else begin
            _T_1280 <= 6'h0;
          end
        end else begin
          _T_1280 <= _T_1282;
        end
      end
    end
    if (reset) begin
      _T_1326 <= 32'h0;
    end else begin
      if (io_in_d_valid) begin
        _T_1326 <= 32'h0;
      end else begin
        _T_1326 <= _T_1337;
      end
    end
    if (reset) begin
      _T_1341 <= 1'h0;
    end else begin
      _T_1341 <= _T_1387;
    end
    if (reset) begin
      _T_1350 <= 6'h0;
    end else begin
      if (io_in_d_valid) begin
        if (_T_1353) begin
          if (_T_1107) begin
            _T_1350 <= _T_1106;
          end else begin
            _T_1350 <= 6'h0;
          end
        end else begin
          _T_1350 <= _T_1352;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel has invalid opcode (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:39 assert (TLMessages.isA(bundle.opcode), \"'A' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:46 assert (visible(edge.address(bundle), bundle.source, edge), \"'A' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:56 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:68 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:77 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:117 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_447) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_447) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_33 & _T_454) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_33 & _T_454) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_33 & _T_458) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_33 & _T_458) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_33 & _T_462) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_33 & _T_462) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_33 & _T_466) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_33 & _T_466) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_33 & _T_470) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_33 & _T_470) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_43 & _T_454) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_43 & _T_454) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_43 & _T_477) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:285 assert (sink_ok, \"'D' channel Grant carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_43 & _T_477) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_43 & _T_458) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_43 & _T_458) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_43 & _T_485) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_43 & _T_485) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_43 & _T_489) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_43 & _T_489) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_43 & _T_466) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_43 & _T_466) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is denied (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:290 assert (deny_put_ok || !bundle.denied, \"'D' channel Grant is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_454) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_55 & _T_454) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_477) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:295 assert (sink_ok, \"'D' channel GrantData carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_55 & _T_477) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_458) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_55 & _T_458) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_485) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_55 & _T_485) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_489) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_55 & _T_489) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_522) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_55 & _T_522) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:300 assert (deny_get_ok || !bundle.denied, \"'D' channel GrantData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_67 & _T_454) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_67 & _T_454) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_67 & _T_462) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_67 & _T_462) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_67 & _T_466) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_67 & _T_466) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is denied (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:308 assert (deny_put_ok || !bundle.denied, \"'D' channel AccessAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_73 & _T_454) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_73 & _T_454) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_73 & _T_462) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_73 & _T_462) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_73 & _T_522) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_73 & _T_522) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:316 assert (deny_get_ok || !bundle.denied, \"'D' channel AccessAckData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_79 & _T_454) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_79 & _T_454) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_79 & _T_462) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_79 & _T_462) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_79 & _T_466) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_79 & _T_466) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is denied (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:324 assert (deny_put_ok || !bundle.denied, \"'D' channel HintAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel has invalid opcode (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:122 assert (TLMessages.isB(bundle.opcode), \"'B' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:124 assert (visible(edge.address(bundle), bundle.source, edge), \"'B' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Probe type unsupported by client (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:133 assert (edge.client.supportsProbe(bundle.source, bundle.size), \"'B' channel carries Probe type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:134 assert (address_ok, \"'B' channel Probe carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries source that is not first source (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:135 assert (legal_source, \"'B' channel Probe carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:136 assert (is_aligned, \"'B' channel Probe address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:137 assert (TLPermissions.isCap(bundle.param), \"'B' channel Probe carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe contains invalid mask (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:138 assert (bundle.mask === mask, \"'B' channel Probe contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe is corrupt (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:139 assert (!bundle.corrupt, \"'B' channel Probe is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Get type unsupported by client (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:143 assert (edge.client.supportsGet(bundle.source, bundle.size), \"'B' channel carries Get type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries unmanaged address (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:144 assert (address_ok, \"'B' channel Get carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries source that is not first source (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:145 assert (legal_source, \"'B' channel Get carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:146 assert (is_aligned, \"'B' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries invalid param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:147 assert (bundle.param === UInt(0), \"'B' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get contains invalid mask (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:148 assert (bundle.mask === mask, \"'B' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get is corrupt (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:149 assert (!bundle.corrupt, \"'B' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutFull type unsupported by client (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:153 assert (edge.client.supportsPutFull(bundle.source, bundle.size), \"'B' channel carries PutFull type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries unmanaged address (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:154 assert (address_ok, \"'B' channel PutFull carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries source that is not first source (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:155 assert (legal_source, \"'B' channel PutFull carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:156 assert (is_aligned, \"'B' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries invalid param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:157 assert (bundle.param === UInt(0), \"'B' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull contains invalid mask (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:158 assert (bundle.mask === mask, \"'B' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutPartial type unsupported by client (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:162 assert (edge.client.supportsPutPartial(bundle.source, bundle.size), \"'B' channel carries PutPartial type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:163 assert (address_ok, \"'B' channel PutPartial carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:164 assert (legal_source, \"'B' channel PutPartial carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:165 assert (is_aligned, \"'B' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries invalid param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:166 assert (bundle.param === UInt(0), \"'B' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial contains invalid mask (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:167 assert ((bundle.mask & ~mask) === UInt(0), \"'B' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Arithmetic type unsupported by client (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:171 assert (edge.client.supportsArithmetic(bundle.source, bundle.size), \"'B' channel carries Arithmetic type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:172 assert (address_ok, \"'B' channel Arithmetic carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:173 assert (legal_source, \"'B' channel Arithmetic carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:174 assert (is_aligned, \"'B' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries invalid opcode param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:175 assert (TLAtomics.isArithmetic(bundle.param), \"'B' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:176 assert (bundle.mask === mask, \"'B' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Logical type unsupported by client (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:180 assert (edge.client.supportsLogical(bundle.source, bundle.size), \"'B' channel carries Logical type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries unmanaged address (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:181 assert (address_ok, \"'B' channel Logical carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries source that is not first source (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:182 assert (legal_source, \"'B' channel Logical carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:183 assert (is_aligned, \"'B' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries invalid opcode param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:184 assert (TLAtomics.isLogical(bundle.param), \"'B' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical contains invalid mask (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:185 assert (bundle.mask === mask, \"'B' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Hint type unsupported by client (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:189 assert (edge.client.supportsHint(bundle.source, bundle.size), \"'B' channel carries Hint type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries unmanaged address (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:190 assert (address_ok, \"'B' channel Hint carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries source that is not first source (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:191 assert (legal_source, \"'B' channel Hint carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:192 assert (is_aligned, \"'B' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint contains invalid mask (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:193 assert (bundle.mask === mask, \"'B' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint is corrupt (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:194 assert (!bundle.corrupt, \"'B' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel has invalid opcode (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:199 assert (TLMessages.isC(bundle.opcode), \"'C' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:205 assert (visible(edge.address(bundle), bundle.source, edge), \"'C' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:208 assert (address_ok, \"'C' channel ProbeAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:209 assert (source_ok, \"'C' channel ProbeAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:210 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:211 assert (is_aligned, \"'C' channel ProbeAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:212 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAck carries invalid report param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck is corrupt (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:213 assert (!bundle.corrupt, \"'C' channel ProbeAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:217 assert (address_ok, \"'C' channel ProbeAckData carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:218 assert (source_ok, \"'C' channel ProbeAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:219 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAckData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:220 assert (is_aligned, \"'C' channel ProbeAckData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:221 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAckData carries invalid report param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:225 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries Release type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:226 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:227 assert (source_ok, \"'C' channel Release carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:228 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel Release smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:229 assert (is_aligned, \"'C' channel Release address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid shrink param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:230 assert (TLPermissions.isShrink(bundle.param), \"'C' channel Release carries invalid shrink param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release is corrupt (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:231 assert (!bundle.corrupt, \"'C' channel Release is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:235 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries ReleaseData type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:236 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:237 assert (source_ok, \"'C' channel ReleaseData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:238 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ReleaseData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:239 assert (is_aligned, \"'C' channel ReleaseData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid shrink param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:240 assert (TLPermissions.isShrink(bundle.param), \"'C' channel ReleaseData carries invalid shrink param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:244 assert (address_ok, \"'C' channel AccessAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:245 assert (source_ok, \"'C' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:246 assert (is_aligned, \"'C' channel AccessAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:247 assert (bundle.param === UInt(0), \"'C' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck is corrupt (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:248 assert (!bundle.corrupt, \"'C' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:252 assert (address_ok, \"'C' channel AccessAckData carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:253 assert (source_ok, \"'C' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:254 assert (is_aligned, \"'C' channel AccessAckData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:255 assert (bundle.param === UInt(0), \"'C' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:259 assert (address_ok, \"'C' channel HintAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:260 assert (source_ok, \"'C' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:261 assert (is_aligned, \"'C' channel HintAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:262 assert (bundle.param === UInt(0), \"'C' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck is corrupt (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:263 assert (!bundle.corrupt, \"'C' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channels carries invalid sink ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:330 assert (sink_ok, \"'E' channels carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1127 & _T_1131) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1127 & _T_1131) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1127 & _T_1135) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1127 & _T_1135) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1127 & _T_1139) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1127 & _T_1139) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1127 & _T_1143) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1127 & _T_1143) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1127 & _T_1147) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1127 & _T_1147) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1127 & _T_1151) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1127 & _T_1151) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel opcode changed within multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:378 assert (b.bits.opcode === opcode, \"'B' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:379 assert (b.bits.param  === param,  \"'B' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel size changed within multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:380 assert (b.bits.size   === size,   \"'B' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel source changed within multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:381 assert (b.bits.source === source, \"'B' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:382 assert (b.bits.address=== address,\"'B' channel addresss changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:401 assert (c.bits.opcode === opcode, \"'C' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:402 assert (c.bits.param  === param,  \"'C' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:403 assert (c.bits.size   === size,   \"'C' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:404 assert (c.bits.source === source, \"'C' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:405 assert (c.bits.address=== address,\"'C' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1308 & _T_1315) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1308 & _T_1315) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1335) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:479 assert (!inflight.orR || limit === UInt(0) || watchdog < limit, \"TileLink timeout expired\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1335) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1368 & _T_1375) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:494 assert(!inflight(bundle.d.bits.sink), \"'D' channel re-used a sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1368 & _T_1375) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at dual_ChipLink.scala:77:31)\n    at Monitor.scala:500 assert((d_set | inflight)(bundle.e.bits.sink), \"'E' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLMonitor_8( 
  input         clock, 
  input         reset, 
  input         io_in_a_ready, 
  input         io_in_a_valid, 
  input  [2:0]  io_in_a_bits_opcode, 
  input  [2:0]  io_in_a_bits_param, 
  input  [2:0]  io_in_a_bits_size, 
  input  [2:0]  io_in_a_bits_source, 
  input  [31:0] io_in_a_bits_address, 
  input  [3:0]  io_in_a_bits_mask, 
  input         io_in_a_bits_corrupt, 
  input         io_in_bvalid, 
  input         io_in_d_ready, 
  input         io_in_d_valid, 
  input  [2:0]  io_in_d_bits_opcode, 
  input  [1:0]  io_in_d_bits_param, 
  input  [2:0]  io_in_d_bits_size, 
  input  [2:0]  io_in_d_bits_source, 
  input  [4:0]  io_in_d_bits_sink, 
  input         io_in_d_bits_denied, 
  input         io_in_d_bits_corrupt 
);
  wire [31:0] plusarg_reader_out; 
  wire  _T_7; 
  wire  _T_8; 
  wire  _T_22; 
  wire [12:0] _T_24; 
  wire [5:0] _T_25; 
  wire [5:0] _T_26; 
  wire [31:0] _GEN_18; 
  wire [31:0] _T_27; 
  wire  _T_28; 
  wire  _T_30; 
  wire [1:0] _T_31; 
  wire [1:0] _T_33; 
  wire  _T_34; 
  wire  _T_35; 
  wire  _T_36; 
  wire  _T_37; 
  wire  _T_39; 
  wire  _T_40; 
  wire  _T_42; 
  wire  _T_43; 
  wire  _T_44; 
  wire  _T_45; 
  wire  _T_46; 
  wire  _T_47; 
  wire  _T_48; 
  wire  _T_49; 
  wire  _T_50; 
  wire  _T_51; 
  wire  _T_52; 
  wire  _T_53; 
  wire  _T_54; 
  wire  _T_55; 
  wire  _T_56; 
  wire  _T_57; 
  wire  _T_58; 
  wire [3:0] _T_61; 
  wire  _T_96; 
  wire [31:0] _T_98; 
  wire [32:0] _T_99; 
  wire [32:0] _T_100; 
  wire [32:0] _T_101; 
  wire  _T_102; 
  wire  _T_104; 
  wire [31:0] _T_106; 
  wire [32:0] _T_107; 
  wire [32:0] _T_108; 
  wire [32:0] _T_109; 
  wire  _T_110; 
  wire  _T_111; 
  wire  _T_115; 
  wire  _T_116; 
  wire  _T_119; 
  wire  _T_121; 
  wire  _T_122; 
  wire  _T_125; 
  wire  _T_126; 
  wire  _T_128; 
  wire  _T_129; 
  wire  _T_130; 
  wire  _T_132; 
  wire  _T_133; 
  wire [3:0] _T_134; 
  wire  _T_135; 
  wire  _T_137; 
  wire  _T_138; 
  wire  _T_139; 
  wire  _T_141; 
  wire  _T_142; 
  wire  _T_143; 
  wire  _T_181; 
  wire  _T_183; 
  wire  _T_184; 
  wire  _T_194; 
  wire  _T_196; 
  wire  _T_209; 
  wire  _T_210; 
  wire  _T_213; 
  wire  _T_214; 
  wire  _T_221; 
  wire  _T_223; 
  wire  _T_224; 
  wire  _T_225; 
  wire  _T_227; 
  wire  _T_228; 
  wire  _T_233; 
  wire  _T_268; 
  wire [3:0] _T_299; 
  wire [3:0] _T_300; 
  wire  _T_301; 
  wire  _T_303; 
  wire  _T_304; 
  wire  _T_305; 
  wire  _T_307; 
  wire  _T_321; 
  wire  _T_324; 
  wire  _T_325; 
  wire  _T_332; 
  wire  _T_334; 
  wire  _T_335; 
  wire  _T_340; 
  wire  _T_367; 
  wire  _T_369; 
  wire  _T_370; 
  wire  _T_375; 
  wire  _T_410; 
  wire  _T_412; 
  wire  _T_413; 
  wire  _T_416; 
  wire  _T_417; 
  wire  _T_431; 
  wire  _T_432; 
  wire  _T_433; 
  wire  _T_435; 
  wire  _T_436; 
  wire  _T_437; 
  wire  _T_439; 
  wire  _T_440; 
  wire  _T_441; 
  wire  _T_443; 
  wire  _T_444; 
  wire  _T_445; 
  wire  _T_447; 
  wire  _T_448; 
  wire  _T_449; 
  wire  _T_451; 
  wire  _T_452; 
  wire  _T_453; 
  wire  _T_458; 
  wire  _T_459; 
  wire  _T_464; 
  wire  _T_466; 
  wire  _T_467; 
  wire  _T_468; 
  wire  _T_470; 
  wire  _T_471; 
  wire  _T_481; 
  wire  _T_501; 
  wire  _T_503; 
  wire  _T_504; 
  wire  _T_510; 
  wire  _T_527; 
  wire  _T_545; 
  wire  _T_562; 
  wire  _T_564; 
  wire  _T_565; 
  wire  _T_574; 
  wire [3:0] _T_579; 
  wire  _T_580; 
  wire  _T_581; 
  reg [3:0] _T_583; 
  reg [31:0] _RAND_0;
  wire [3:0] _T_585; 
  wire  _T_586; 
  reg [2:0] _T_594; 
  reg [31:0] _RAND_1;
  reg [2:0] _T_595; 
  reg [31:0] _RAND_2;
  reg [2:0] _T_596; 
  reg [31:0] _RAND_3;
  reg [2:0] _T_597; 
  reg [31:0] _RAND_4;
  reg [31:0] _T_598; 
  reg [31:0] _RAND_5;
  wire  _T_599; 
  wire  _T_600; 
  wire  _T_601; 
  wire  _T_603; 
  wire  _T_604; 
  wire  _T_605; 
  wire  _T_607; 
  wire  _T_608; 
  wire  _T_609; 
  wire  _T_611; 
  wire  _T_612; 
  wire  _T_613; 
  wire  _T_615; 
  wire  _T_616; 
  wire  _T_617; 
  wire  _T_619; 
  wire  _T_620; 
  wire  _T_622; 
  wire  _T_623; 
  wire [12:0] _T_625; 
  wire [5:0] _T_626; 
  wire [5:0] _T_627; 
  wire [3:0] _T_628; 
  wire  _T_629; 
  reg [3:0] _T_631; 
  reg [31:0] _RAND_6;
  wire [3:0] _T_633; 
  wire  _T_634; 
  reg [2:0] _T_642; 
  reg [31:0] _RAND_7;
  reg [1:0] _T_643; 
  reg [31:0] _RAND_8;
  reg [2:0] _T_644; 
  reg [31:0] _RAND_9;
  reg [2:0] _T_645; 
  reg [31:0] _RAND_10;
  reg [4:0] _T_646; 
  reg [31:0] _RAND_11;
  reg  _T_647; 
  reg [31:0] _RAND_12;
  wire  _T_648; 
  wire  _T_649; 
  wire  _T_650; 
  wire  _T_652; 
  wire  _T_653; 
  wire  _T_654; 
  wire  _T_656; 
  wire  _T_657; 
  wire  _T_658; 
  wire  _T_660; 
  wire  _T_661; 
  wire  _T_662; 
  wire  _T_664; 
  wire  _T_665; 
  wire  _T_666; 
  wire  _T_668; 
  wire  _T_669; 
  wire  _T_670; 
  wire  _T_672; 
  wire  _T_673; 
  wire  _T_675; 
  reg [7:0] _T_676; 
  reg [31:0] _RAND_13;
  reg [3:0] _T_686; 
  reg [31:0] _RAND_14;
  wire [3:0] _T_688; 
  wire  _T_689; 
  reg [3:0] _T_705; 
  reg [31:0] _RAND_15;
  wire [3:0] _T_707; 
  wire  _T_708; 
  wire  _T_718; 
  wire [7:0] _T_720; 
  wire [7:0] _T_721; 
  wire  _T_722; 
  wire  _T_723; 
  wire  _T_725; 
  wire  _T_726; 
  wire [7:0] _GEN_15; 
  wire  _T_730; 
  wire  _T_732; 
  wire  _T_733; 
  wire [7:0] _T_734; 
  wire [7:0] _T_735; 
  wire [7:0] _T_736; 
  wire  _T_737; 
  wire  _T_739; 
  wire  _T_740; 
  wire [7:0] _GEN_16; 
  wire  _T_741; 
  wire  _T_742; 
  wire  _T_743; 
  wire  _T_744; 
  wire  _T_746; 
  wire  _T_747; 
  wire [7:0] _T_748; 
  wire [7:0] _T_749; 
  wire [7:0] _T_750; 
  reg [31:0] _T_751; 
  reg [31:0] _RAND_16;
  wire  _T_752; 
  wire  _T_753; 
  wire  _T_754; 
  wire  _T_755; 
  wire  _T_756; 
  wire  _T_757; 
  wire  _T_759; 
  wire  _T_760; 
  wire [31:0] _T_762; 
  wire  _T_765; 
  wire  _GEN_19; 
  wire  _GEN_35; 
  wire  _GEN_53; 
  wire  _GEN_65; 
  wire  _GEN_75; 
  wire  _GEN_85; 
  wire  _GEN_95; 
  wire  _GEN_105; 
  wire  _GEN_115; 
  wire  _GEN_125; 
  wire  _GEN_137; 
  wire  _GEN_149; 
  wire  _GEN_155; 
  wire  _GEN_161; 
  dual_plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0)) plusarg_reader ( 
    .out(plusarg_reader_out)
  );
  assign _T_7 = io_in_a_bits_source[2:2]; 
  assign _T_8 = _T_7 == 1'h0; 
  assign _T_22 = _T_8 | _T_7; 
  assign _T_24 = 13'h3f << io_in_a_bits_size; 
  assign _T_25 = _T_24[5:0]; 
  assign _T_26 = ~ _T_25; 
  assign _GEN_18 = {{26'd0}, _T_26}; 
  assign _T_27 = io_in_a_bits_address & _GEN_18; 
  assign _T_28 = _T_27 == 32'h0; 
  assign _T_30 = io_in_a_bits_size[0]; 
  assign _T_31 = 2'h1 << _T_30; 
  assign _T_33 = _T_31 | 2'h1; 
  assign _T_34 = io_in_a_bits_size >= 3'h2; 
  assign _T_35 = _T_33[1]; 
  assign _T_36 = io_in_a_bits_address[1]; 
  assign _T_37 = _T_36 == 1'h0; 
  assign _T_39 = _T_35 & _T_37; 
  assign _T_40 = _T_34 | _T_39; 
  assign _T_42 = _T_35 & _T_36; 
  assign _T_43 = _T_34 | _T_42; 
  assign _T_44 = _T_33[0]; 
  assign _T_45 = io_in_a_bits_address[0]; 
  assign _T_46 = _T_45 == 1'h0; 
  assign _T_47 = _T_37 & _T_46; 
  assign _T_48 = _T_44 & _T_47; 
  assign _T_49 = _T_40 | _T_48; 
  assign _T_50 = _T_37 & _T_45; 
  assign _T_51 = _T_44 & _T_50; 
  assign _T_52 = _T_40 | _T_51; 
  assign _T_53 = _T_36 & _T_46; 
  assign _T_54 = _T_44 & _T_53; 
  assign _T_55 = _T_43 | _T_54; 
  assign _T_56 = _T_36 & _T_45; 
  assign _T_57 = _T_44 & _T_56; 
  assign _T_58 = _T_43 | _T_57; 
  assign _T_61 = {_T_58,_T_55,_T_52,_T_49}; 
  assign _T_96 = io_in_a_bits_opcode == 3'h6; 
  assign _T_98 = io_in_a_bits_address ^ 32'h40000000; 
  assign _T_99 = {1'b0,$signed(_T_98)}; 
  assign _T_100 = $signed(_T_99) & $signed(-33'sh20000000); 
  assign _T_101 = $signed(_T_100); 
  assign _T_102 = $signed(_T_101) == $signed(33'sh0); 
  assign _T_104 = 3'h6 == io_in_a_bits_size; 
  assign _T_106 = io_in_a_bits_address ^ 32'h80000000; 
  assign _T_107 = {1'b0,$signed(_T_106)}; 
  assign _T_108 = $signed(_T_107) & $signed(-33'sh80000000); 
  assign _T_109 = $signed(_T_108); 
  assign _T_110 = $signed(_T_109) == $signed(33'sh0); 
  assign _T_111 = _T_104 & _T_110; 
  assign _T_115 = _T_111 | reset; 
  assign _T_116 = _T_115 == 1'h0; 
  assign _T_119 = reset == 1'h0; 
  assign _T_121 = _T_22 | reset; 
  assign _T_122 = _T_121 == 1'h0; 
  assign _T_125 = _T_34 | reset; 
  assign _T_126 = _T_125 == 1'h0; 
  assign _T_128 = _T_28 | reset; 
  assign _T_129 = _T_128 == 1'h0; 
  assign _T_130 = io_in_a_bits_param <= 3'h2; 
  assign _T_132 = _T_130 | reset; 
  assign _T_133 = _T_132 == 1'h0; 
  assign _T_134 = ~ io_in_a_bits_mask; 
  assign _T_135 = _T_134 == 4'h0; 
  assign _T_137 = _T_135 | reset; 
  assign _T_138 = _T_137 == 1'h0; 
  assign _T_139 = io_in_a_bits_corrupt == 1'h0; 
  assign _T_141 = _T_139 | reset; 
  assign _T_142 = _T_141 == 1'h0; 
  assign _T_143 = io_in_a_bits_opcode == 3'h7; 
  assign _T_181 = io_in_a_bits_param != 3'h0; 
  assign _T_183 = _T_181 | reset; 
  assign _T_184 = _T_183 == 1'h0; 
  assign _T_194 = io_in_a_bits_opcode == 3'h4; 
  assign _T_196 = io_in_a_bits_size <= 3'h6; 
  assign _T_209 = _T_102 | _T_110; 
  assign _T_210 = _T_196 & _T_209; 
  assign _T_213 = _T_210 | reset; 
  assign _T_214 = _T_213 == 1'h0; 
  assign _T_221 = io_in_a_bits_param == 3'h0; 
  assign _T_223 = _T_221 | reset; 
  assign _T_224 = _T_223 == 1'h0; 
  assign _T_225 = io_in_a_bits_mask == _T_61; 
  assign _T_227 = _T_225 | reset; 
  assign _T_228 = _T_227 == 1'h0; 
  assign _T_233 = io_in_a_bits_opcode == 3'h0; 
  assign _T_268 = io_in_a_bits_opcode == 3'h1; 
  assign _T_299 = ~ _T_61; 
  assign _T_300 = io_in_a_bits_mask & _T_299; 
  assign _T_301 = _T_300 == 4'h0; 
  assign _T_303 = _T_301 | reset; 
  assign _T_304 = _T_303 == 1'h0; 
  assign _T_305 = io_in_a_bits_opcode == 3'h2; 
  assign _T_307 = io_in_a_bits_size <= 3'h3; 
  assign _T_321 = _T_307 & _T_209; 
  assign _T_324 = _T_321 | reset; 
  assign _T_325 = _T_324 == 1'h0; 
  assign _T_332 = io_in_a_bits_param <= 3'h4; 
  assign _T_334 = _T_332 | reset; 
  assign _T_335 = _T_334 == 1'h0; 
  assign _T_340 = io_in_a_bits_opcode == 3'h3; 
  assign _T_367 = io_in_a_bits_param <= 3'h3; 
  assign _T_369 = _T_367 | reset; 
  assign _T_370 = _T_369 == 1'h0; 
  assign _T_375 = io_in_a_bits_opcode == 3'h5; 
  assign _T_410 = io_in_d_bits_opcode <= 3'h6; 
  assign _T_412 = _T_410 | reset; 
  assign _T_413 = _T_412 == 1'h0; 
  assign _T_416 = io_in_d_bits_source[2:2]; 
  assign _T_417 = _T_416 == 1'h0; 
  assign _T_431 = _T_417 | _T_416; 
  assign _T_432 = io_in_d_bits_sink < 5'h1f; 
  assign _T_433 = io_in_d_bits_opcode == 3'h6; 
  assign _T_435 = _T_431 | reset; 
  assign _T_436 = _T_435 == 1'h0; 
  assign _T_437 = io_in_d_bits_size >= 3'h2; 
  assign _T_439 = _T_437 | reset; 
  assign _T_440 = _T_439 == 1'h0; 
  assign _T_441 = io_in_d_bits_param == 2'h0; 
  assign _T_443 = _T_441 | reset; 
  assign _T_444 = _T_443 == 1'h0; 
  assign _T_445 = io_in_d_bits_corrupt == 1'h0; 
  assign _T_447 = _T_445 | reset; 
  assign _T_448 = _T_447 == 1'h0; 
  assign _T_449 = io_in_d_bits_denied == 1'h0; 
  assign _T_451 = _T_449 | reset; 
  assign _T_452 = _T_451 == 1'h0; 
  assign _T_453 = io_in_d_bits_opcode == 3'h4; 
  assign _T_458 = _T_432 | reset; 
  assign _T_459 = _T_458 == 1'h0; 
  assign _T_464 = io_in_d_bits_param <= 2'h2; 
  assign _T_466 = _T_464 | reset; 
  assign _T_467 = _T_466 == 1'h0; 
  assign _T_468 = io_in_d_bits_param != 2'h2; 
  assign _T_470 = _T_468 | reset; 
  assign _T_471 = _T_470 == 1'h0; 
  assign _T_481 = io_in_d_bits_opcode == 3'h5; 
  assign _T_501 = _T_449 | io_in_d_bits_corrupt; 
  assign _T_503 = _T_501 | reset; 
  assign _T_504 = _T_503 == 1'h0; 
  assign _T_510 = io_in_d_bits_opcode == 3'h0; 
  assign _T_527 = io_in_d_bits_opcode == 3'h1; 
  assign _T_545 = io_in_d_bits_opcode == 3'h2; 
  assign _T_562 = io_in_bvalid == 1'h0; 
  assign _T_564 = _T_562 | reset; 
  assign _T_565 = _T_564 == 1'h0; 
  assign _T_574 = io_in_a_ready & io_in_a_valid; 
  assign _T_579 = _T_26[5:2]; 
  assign _T_580 = io_in_a_bits_opcode[2]; 
  assign _T_581 = _T_580 == 1'h0; 
  assign _T_585 = _T_583 - 4'h1; 
  assign _T_586 = _T_583 == 4'h0; 
  assign _T_599 = _T_586 == 1'h0; 
  assign _T_600 = io_in_a_valid & _T_599; 
  assign _T_601 = io_in_a_bits_opcode == _T_594; 
  assign _T_603 = _T_601 | reset; 
  assign _T_604 = _T_603 == 1'h0; 
  assign _T_605 = io_in_a_bits_param == _T_595; 
  assign _T_607 = _T_605 | reset; 
  assign _T_608 = _T_607 == 1'h0; 
  assign _T_609 = io_in_a_bits_size == _T_596; 
  assign _T_611 = _T_609 | reset; 
  assign _T_612 = _T_611 == 1'h0; 
  assign _T_613 = io_in_a_bits_source == _T_597; 
  assign _T_615 = _T_613 | reset; 
  assign _T_616 = _T_615 == 1'h0; 
  assign _T_617 = io_in_a_bits_address == _T_598; 
  assign _T_619 = _T_617 | reset; 
  assign _T_620 = _T_619 == 1'h0; 
  assign _T_622 = _T_574 & _T_586; 
  assign _T_623 = io_in_d_ready & io_in_d_valid; 
  assign _T_625 = 13'h3f << io_in_d_bits_size; 
  assign _T_626 = _T_625[5:0]; 
  assign _T_627 = ~ _T_626; 
  assign _T_628 = _T_627[5:2]; 
  assign _T_629 = io_in_d_bits_opcode[0]; 
  assign _T_633 = _T_631 - 4'h1; 
  assign _T_634 = _T_631 == 4'h0; 
  assign _T_648 = _T_634 == 1'h0; 
  assign _T_649 = io_in_d_valid & _T_648; 
  assign _T_650 = io_in_d_bits_opcode == _T_642; 
  assign _T_652 = _T_650 | reset; 
  assign _T_653 = _T_652 == 1'h0; 
  assign _T_654 = io_in_d_bits_param == _T_643; 
  assign _T_656 = _T_654 | reset; 
  assign _T_657 = _T_656 == 1'h0; 
  assign _T_658 = io_in_d_bits_size == _T_644; 
  assign _T_660 = _T_658 | reset; 
  assign _T_661 = _T_660 == 1'h0; 
  assign _T_662 = io_in_d_bits_source == _T_645; 
  assign _T_664 = _T_662 | reset; 
  assign _T_665 = _T_664 == 1'h0; 
  assign _T_666 = io_in_d_bits_sink == _T_646; 
  assign _T_668 = _T_666 | reset; 
  assign _T_669 = _T_668 == 1'h0; 
  assign _T_670 = io_in_d_bits_denied == _T_647; 
  assign _T_672 = _T_670 | reset; 
  assign _T_673 = _T_672 == 1'h0; 
  assign _T_675 = _T_623 & _T_634; 
  assign _T_688 = _T_686 - 4'h1; 
  assign _T_689 = _T_686 == 4'h0; 
  assign _T_707 = _T_705 - 4'h1; 
  assign _T_708 = _T_705 == 4'h0; 
  assign _T_718 = _T_574 & _T_689; 
  assign _T_720 = 8'h1 << io_in_a_bits_source; 
  assign _T_721 = _T_676 >> io_in_a_bits_source; 
  assign _T_722 = _T_721[0]; 
  assign _T_723 = _T_722 == 1'h0; 
  assign _T_725 = _T_723 | reset; 
  assign _T_726 = _T_725 == 1'h0; 
  assign _GEN_15 = _T_718 ? _T_720 : 8'h0; 
  assign _T_730 = _T_623 & _T_708; 
  assign _T_732 = _T_433 == 1'h0; 
  assign _T_733 = _T_730 & _T_732; 
  assign _T_734 = 8'h1 << io_in_d_bits_source; 
  assign _T_735 = _GEN_15 | _T_676; 
  assign _T_736 = _T_735 >> io_in_d_bits_source; 
  assign _T_737 = _T_736[0]; 
  assign _T_739 = _T_737 | reset; 
  assign _T_740 = _T_739 == 1'h0; 
  assign _GEN_16 = _T_733 ? _T_734 : 8'h0; 
  assign _T_741 = _GEN_15 != _GEN_16; 
  assign _T_742 = _GEN_15 != 8'h0; 
  assign _T_743 = _T_742 == 1'h0; 
  assign _T_744 = _T_741 | _T_743; 
  assign _T_746 = _T_744 | reset; 
  assign _T_747 = _T_746 == 1'h0; 
  assign _T_748 = _T_676 | _GEN_15; 
  assign _T_749 = ~ _GEN_16; 
  assign _T_750 = _T_748 & _T_749; 
  assign _T_752 = _T_676 != 8'h0; 
  assign _T_753 = _T_752 == 1'h0; 
  assign _T_754 = plusarg_reader_out == 32'h0; 
  assign _T_755 = _T_753 | _T_754; 
  assign _T_756 = _T_751 < plusarg_reader_out; 
  assign _T_757 = _T_755 | _T_756; 
  assign _T_759 = _T_757 | reset; 
  assign _T_760 = _T_759 == 1'h0; 
  assign _T_762 = _T_751 + 32'h1; 
  assign _T_765 = _T_574 | _T_623; 
  assign _GEN_19 = io_in_a_valid & _T_96; 
  assign _GEN_35 = io_in_a_valid & _T_143; 
  assign _GEN_53 = io_in_a_valid & _T_194; 
  assign _GEN_65 = io_in_a_valid & _T_233; 
  assign _GEN_75 = io_in_a_valid & _T_268; 
  assign _GEN_85 = io_in_a_valid & _T_305; 
  assign _GEN_95 = io_in_a_valid & _T_340; 
  assign _GEN_105 = io_in_a_valid & _T_375; 
  assign _GEN_115 = io_in_d_valid & _T_433; 
  assign _GEN_125 = io_in_d_valid & _T_453; 
  assign _GEN_137 = io_in_d_valid & _T_481; 
  assign _GEN_149 = io_in_d_valid & _T_510; 
  assign _GEN_155 = io_in_d_valid & _T_527; 
  assign _GEN_161 = io_in_d_valid & _T_545; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_583 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_594 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_595 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_596 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_597 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_598 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_631 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_642 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_643 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_644 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_645 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_646 = _RAND_11[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_647 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_676 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_686 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_705 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_751 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_583 <= 4'h0;
    end else begin
      if (_T_574) begin
        if (_T_586) begin
          if (_T_581) begin
            _T_583 <= _T_579;
          end else begin
            _T_583 <= 4'h0;
          end
        end else begin
          _T_583 <= _T_585;
        end
      end
    end
    if (_T_622) begin
      _T_594 <= io_in_a_bits_opcode;
    end
    if (_T_622) begin
      _T_595 <= io_in_a_bits_param;
    end
    if (_T_622) begin
      _T_596 <= io_in_a_bits_size;
    end
    if (_T_622) begin
      _T_597 <= io_in_a_bits_source;
    end
    if (_T_622) begin
      _T_598 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_631 <= 4'h0;
    end else begin
      if (_T_623) begin
        if (_T_634) begin
          if (_T_629) begin
            _T_631 <= _T_628;
          end else begin
            _T_631 <= 4'h0;
          end
        end else begin
          _T_631 <= _T_633;
        end
      end
    end
    if (_T_675) begin
      _T_642 <= io_in_d_bits_opcode;
    end
    if (_T_675) begin
      _T_643 <= io_in_d_bits_param;
    end
    if (_T_675) begin
      _T_644 <= io_in_d_bits_size;
    end
    if (_T_675) begin
      _T_645 <= io_in_d_bits_source;
    end
    if (_T_675) begin
      _T_646 <= io_in_d_bits_sink;
    end
    if (_T_675) begin
      _T_647 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_676 <= 8'h0;
    end else begin
      _T_676 <= _T_750;
    end
    if (reset) begin
      _T_686 <= 4'h0;
    end else begin
      if (_T_574) begin
        if (_T_689) begin
          if (_T_581) begin
            _T_686 <= _T_579;
          end else begin
            _T_686 <= 4'h0;
          end
        end else begin
          _T_686 <= _T_688;
        end
      end
    end
    if (reset) begin
      _T_705 <= 4'h0;
    end else begin
      if (_T_623) begin
        if (_T_708) begin
          if (_T_629) begin
            _T_705 <= _T_628;
          end else begin
            _T_705 <= 4'h0;
          end
        end else begin
          _T_705 <= _T_707;
        end
      end
    end
    if (reset) begin
      _T_751 <= 32'h0;
    end else begin
      if (_T_765) begin
        _T_751 <= 32'h0;
      end else begin
        _T_751 <= _T_762;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel has invalid opcode (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:39 assert (TLMessages.isA(bundle.opcode), \"'A' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:46 assert (visible(edge.address(bundle), bundle.source, edge), \"'A' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_119) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_119) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_122) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_122) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_126) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_126) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_129) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_138) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_138) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_142) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:56 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_142) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_116) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_119) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_119) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_122) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_122) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_126) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_126) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_129) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_133) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_184) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_184) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_138) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_138) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_142) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:68 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_142) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_214) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_214) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_122) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_122) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_129) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_224) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_224) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_228) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_228) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_142) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:77 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_142) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_214) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_214) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_122) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_122) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_129) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_224) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_224) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_228) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_228) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_214) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_214) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_122) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_122) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_129) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_224) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_224) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_304) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_304) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_325) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_325) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_122) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_122) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_129) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_335) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_335) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_228) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_228) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_325) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_325) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_122) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_122) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_129) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_370) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_370) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_228) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_228) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_214) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_214) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_122) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_122) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_129) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_228) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_228) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_142) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:117 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_142) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_413) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_413) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_436) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_436) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_440) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_440) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_444) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_444) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_448) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_448) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_452) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_452) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_436) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_436) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_459) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:285 assert (sink_ok, \"'D' channel Grant carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_459) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_440) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_440) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_467) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_467) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_471) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_471) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & _T_448) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & _T_448) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is denied (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:290 assert (deny_put_ok || !bundle.denied, \"'D' channel Grant is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_436) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_436) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_459) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:295 assert (sink_ok, \"'D' channel GrantData carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_459) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_440) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_440) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_467) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_467) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_471) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_471) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_137 & _T_504) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_137 & _T_504) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:300 assert (deny_get_ok || !bundle.denied, \"'D' channel GrantData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_436) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_436) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_444) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_444) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_149 & _T_448) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_149 & _T_448) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is denied (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:308 assert (deny_put_ok || !bundle.denied, \"'D' channel AccessAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_436) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_436) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_444) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_444) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_155 & _T_504) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_155 & _T_504) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:316 assert (deny_get_ok || !bundle.denied, \"'D' channel AccessAckData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_436) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_436) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_444) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_444) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_448) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_448) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is denied (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:324 assert (deny_put_ok || !bundle.denied, \"'D' channel HintAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_565) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel valid and not TL-C (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:341 assert (!bundle.b.valid, \"'B' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_565) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel valid and not TL-C (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:342 assert (!bundle.c.valid, \"'C' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel valid and not TL-C (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:343 assert (!bundle.e.valid, \"'E' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_600 & _T_604) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_600 & _T_604) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_600 & _T_608) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_600 & _T_608) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_600 & _T_612) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_600 & _T_612) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_600 & _T_616) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_600 & _T_616) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_600 & _T_620) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_600 & _T_620) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_649 & _T_653) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_649 & _T_653) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_649 & _T_657) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_649 & _T_657) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_649 & _T_661) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_649 & _T_661) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_649 & _T_665) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_649 & _T_665) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_649 & _T_669) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_649 & _T_669) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_649 & _T_673) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_649 & _T_673) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_718 & _T_726) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_718 & _T_726) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_733 & _T_740) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_733 & _T_740) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_747) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 8 (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_747) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_760) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at dual_ChipLink.scala:67:13)\n    at Monitor.scala:479 assert (!inflight.orR || limit === UInt(0) || watchdog < limit, \"TileLink timeout expired\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_760) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLMonitor_9( 
  input         clock, 
  input         reset, 
  input         io_in_a_ready, 
  input         io_in_a_valid, 
  input  [2:0]  io_in_a_bits_opcode, 
  input  [2:0]  io_in_a_bits_param, 
  input  [2:0]  io_in_a_bits_size, 
  input  [6:0]  io_in_a_bits_source, 
  input  [31:0] io_in_a_bits_address, 
  input  [7:0]  io_in_a_bits_mask, 
  input         io_in_a_bits_corrupt, 
  input         io_in_d_ready, 
  input         io_in_d_valid, 
  input  [2:0]  io_in_d_bits_opcode, 
  input  [2:0]  io_in_d_bits_size, 
  input  [6:0]  io_in_d_bits_source, 
  input         io_in_d_bits_denied, 
  input         io_in_d_bits_corrupt 
);
  wire [31:0] plusarg_reader_out; 
  wire [2:0] _T_7; 
  wire  _T_8; 
  wire  _T_16; 
  wire  _T_24; 
  wire  _T_32; 
  wire  _T_40; 
  wire  _T_48; 
  wire  _T_56; 
  wire  _T_64; 
  wire  _T_70; 
  wire  _T_71; 
  wire  _T_72; 
  wire  _T_73; 
  wire  _T_74; 
  wire  _T_75; 
  wire  _T_76; 
  wire [12:0] _T_78; 
  wire [5:0] _T_79; 
  wire [5:0] _T_80; 
  wire [31:0] _GEN_18; 
  wire [31:0] _T_81; 
  wire  _T_82; 
  wire [1:0] _T_84; 
  wire [3:0] _T_85; 
  wire [2:0] _T_86; 
  wire [2:0] _T_87; 
  wire  _T_88; 
  wire  _T_89; 
  wire  _T_90; 
  wire  _T_91; 
  wire  _T_93; 
  wire  _T_94; 
  wire  _T_96; 
  wire  _T_97; 
  wire  _T_98; 
  wire  _T_99; 
  wire  _T_100; 
  wire  _T_101; 
  wire  _T_102; 
  wire  _T_103; 
  wire  _T_104; 
  wire  _T_105; 
  wire  _T_106; 
  wire  _T_107; 
  wire  _T_108; 
  wire  _T_109; 
  wire  _T_110; 
  wire  _T_111; 
  wire  _T_112; 
  wire  _T_113; 
  wire  _T_114; 
  wire  _T_115; 
  wire  _T_116; 
  wire  _T_117; 
  wire  _T_118; 
  wire  _T_119; 
  wire  _T_120; 
  wire  _T_121; 
  wire  _T_122; 
  wire  _T_123; 
  wire  _T_124; 
  wire  _T_125; 
  wire  _T_126; 
  wire  _T_127; 
  wire  _T_128; 
  wire  _T_129; 
  wire  _T_130; 
  wire  _T_131; 
  wire  _T_132; 
  wire  _T_133; 
  wire  _T_134; 
  wire  _T_135; 
  wire  _T_136; 
  wire  _T_137; 
  wire  _T_138; 
  wire  _T_139; 
  wire [7:0] _T_146; 
  wire  _T_277; 
  wire [31:0] _T_279; 
  wire [32:0] _T_280; 
  wire [32:0] _T_281; 
  wire [32:0] _T_282; 
  wire  _T_283; 
  wire  _T_288; 
  wire  _T_355; 
  wire  _T_357; 
  wire  _T_374; 
  wire  _T_375; 
  wire  _T_377; 
  wire  _T_378; 
  wire  _T_381; 
  wire  _T_382; 
  wire  _T_384; 
  wire  _T_385; 
  wire  _T_386; 
  wire  _T_388; 
  wire  _T_389; 
  wire [7:0] _T_390; 
  wire  _T_391; 
  wire  _T_393; 
  wire  _T_394; 
  wire  _T_395; 
  wire  _T_397; 
  wire  _T_398; 
  wire  _T_399; 
  wire  _T_512; 
  wire  _T_514; 
  wire  _T_515; 
  wire  _T_525; 
  wire  _T_535; 
  wire  _T_538; 
  wire  _T_539; 
  wire  _T_546; 
  wire  _T_548; 
  wire  _T_549; 
  wire  _T_550; 
  wire  _T_552; 
  wire  _T_553; 
  wire  _T_558; 
  wire  _T_587; 
  wire [7:0] _T_612; 
  wire [7:0] _T_613; 
  wire  _T_614; 
  wire  _T_616; 
  wire  _T_617; 
  wire  _T_618; 
  wire  _T_636; 
  wire  _T_638; 
  wire  _T_639; 
  wire  _T_644; 
  wire  _T_662; 
  wire  _T_664; 
  wire  _T_665; 
  wire  _T_670; 
  wire  _T_696; 
  wire  _T_698; 
  wire  _T_699; 
  wire [2:0] _T_702; 
  wire  _T_703; 
  wire  _T_711; 
  wire  _T_719; 
  wire  _T_727; 
  wire  _T_735; 
  wire  _T_743; 
  wire  _T_751; 
  wire  _T_759; 
  wire  _T_765; 
  wire  _T_766; 
  wire  _T_767; 
  wire  _T_768; 
  wire  _T_769; 
  wire  _T_770; 
  wire  _T_771; 
  wire  _T_773; 
  wire  _T_775; 
  wire  _T_776; 
  wire  _T_777; 
  wire  _T_779; 
  wire  _T_780; 
  wire  _T_785; 
  wire  _T_787; 
  wire  _T_788; 
  wire  _T_789; 
  wire  _T_791; 
  wire  _T_792; 
  wire  _T_793; 
  wire  _T_821; 
  wire  _T_841; 
  wire  _T_843; 
  wire  _T_844; 
  wire  _T_850; 
  wire  _T_867; 
  wire  _T_885; 
  wire  _T_914; 
  wire [2:0] _T_919; 
  wire  _T_920; 
  wire  _T_921; 
  reg [2:0] _T_923; 
  reg [31:0] _RAND_0;
  wire [2:0] _T_925; 
  wire  _T_926; 
  reg [2:0] _T_934; 
  reg [31:0] _RAND_1;
  reg [2:0] _T_935; 
  reg [31:0] _RAND_2;
  reg [2:0] _T_936; 
  reg [31:0] _RAND_3;
  reg [6:0] _T_937; 
  reg [31:0] _RAND_4;
  reg [31:0] _T_938; 
  reg [31:0] _RAND_5;
  wire  _T_939; 
  wire  _T_940; 
  wire  _T_941; 
  wire  _T_943; 
  wire  _T_944; 
  wire  _T_945; 
  wire  _T_947; 
  wire  _T_948; 
  wire  _T_949; 
  wire  _T_951; 
  wire  _T_952; 
  wire  _T_953; 
  wire  _T_955; 
  wire  _T_956; 
  wire  _T_957; 
  wire  _T_959; 
  wire  _T_960; 
  wire  _T_962; 
  wire  _T_963; 
  wire [12:0] _T_965; 
  wire [5:0] _T_966; 
  wire [5:0] _T_967; 
  wire [2:0] _T_968; 
  wire  _T_969; 
  reg [2:0] _T_971; 
  reg [31:0] _RAND_6;
  wire [2:0] _T_973; 
  wire  _T_974; 
  reg [2:0] _T_982; 
  reg [31:0] _RAND_7;
  reg [2:0] _T_984; 
  reg [31:0] _RAND_8;
  reg [6:0] _T_985; 
  reg [31:0] _RAND_9;
  reg  _T_987; 
  reg [31:0] _RAND_10;
  wire  _T_988; 
  wire  _T_989; 
  wire  _T_990; 
  wire  _T_992; 
  wire  _T_993; 
  wire  _T_998; 
  wire  _T_1000; 
  wire  _T_1001; 
  wire  _T_1002; 
  wire  _T_1004; 
  wire  _T_1005; 
  wire  _T_1010; 
  wire  _T_1012; 
  wire  _T_1013; 
  wire  _T_1015; 
  reg [127:0] _T_1016; 
  reg [127:0] _RAND_11;
  reg [2:0] _T_1026; 
  reg [31:0] _RAND_12;
  wire [2:0] _T_1028; 
  wire  _T_1029; 
  reg [2:0] _T_1045; 
  reg [31:0] _RAND_13;
  wire [2:0] _T_1047; 
  wire  _T_1048; 
  wire  _T_1058; 
  wire [127:0] _T_1060; 
  wire [127:0] _T_1061; 
  wire  _T_1062; 
  wire  _T_1063; 
  wire  _T_1065; 
  wire  _T_1066; 
  wire [127:0] _GEN_15; 
  wire  _T_1070; 
  wire  _T_1072; 
  wire  _T_1073; 
  wire [127:0] _T_1074; 
  wire [127:0] _T_1075; 
  wire [127:0] _T_1076; 
  wire  _T_1077; 
  wire  _T_1079; 
  wire  _T_1080; 
  wire [127:0] _GEN_16; 
  wire  _T_1081; 
  wire  _T_1082; 
  wire  _T_1083; 
  wire  _T_1084; 
  wire  _T_1086; 
  wire  _T_1087; 
  wire [127:0] _T_1088; 
  wire [127:0] _T_1089; 
  wire [127:0] _T_1090; 
  reg [31:0] _T_1091; 
  reg [31:0] _RAND_14;
  wire  _T_1092; 
  wire  _T_1093; 
  wire  _T_1094; 
  wire  _T_1095; 
  wire  _T_1096; 
  wire  _T_1097; 
  wire  _T_1099; 
  wire  _T_1100; 
  wire [31:0] _T_1102; 
  wire  _T_1105; 
  wire  _GEN_19; 
  wire  _GEN_35; 
  wire  _GEN_53; 
  wire  _GEN_65; 
  wire  _GEN_75; 
  wire  _GEN_85; 
  wire  _GEN_95; 
  wire  _GEN_105; 
  wire  _GEN_115; 
  wire  _GEN_123; 
  wire  _GEN_131; 
  wire  _GEN_139; 
  wire  _GEN_143; 
  wire  _GEN_147; 
  dual_plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0)) plusarg_reader ( 
    .out(plusarg_reader_out)
  );
  assign _T_7 = io_in_a_bits_source[6:4]; 
  assign _T_8 = _T_7 == 3'h0; 
  assign _T_16 = _T_7 == 3'h1; 
  assign _T_24 = _T_7 == 3'h2; 
  assign _T_32 = _T_7 == 3'h3; 
  assign _T_40 = _T_7 == 3'h4; 
  assign _T_48 = _T_7 == 3'h5; 
  assign _T_56 = _T_7 == 3'h6; 
  assign _T_64 = _T_7 == 3'h7; 
  assign _T_70 = _T_8 | _T_16; 
  assign _T_71 = _T_70 | _T_24; 
  assign _T_72 = _T_71 | _T_32; 
  assign _T_73 = _T_72 | _T_40; 
  assign _T_74 = _T_73 | _T_48; 
  assign _T_75 = _T_74 | _T_56; 
  assign _T_76 = _T_75 | _T_64; 
  assign _T_78 = 13'h3f << io_in_a_bits_size; 
  assign _T_79 = _T_78[5:0]; 
  assign _T_80 = ~ _T_79; 
  assign _GEN_18 = {{26'd0}, _T_80}; 
  assign _T_81 = io_in_a_bits_address & _GEN_18; 
  assign _T_82 = _T_81 == 32'h0; 
  assign _T_84 = io_in_a_bits_size[1:0]; 
  assign _T_85 = 4'h1 << _T_84; 
  assign _T_86 = _T_85[2:0]; 
  assign _T_87 = _T_86 | 3'h1; 
  assign _T_88 = io_in_a_bits_size >= 3'h3; 
  assign _T_89 = _T_87[2]; 
  assign _T_90 = io_in_a_bits_address[2]; 
  assign _T_91 = _T_90 == 1'h0; 
  assign _T_93 = _T_89 & _T_91; 
  assign _T_94 = _T_88 | _T_93; 
  assign _T_96 = _T_89 & _T_90; 
  assign _T_97 = _T_88 | _T_96; 
  assign _T_98 = _T_87[1]; 
  assign _T_99 = io_in_a_bits_address[1]; 
  assign _T_100 = _T_99 == 1'h0; 
  assign _T_101 = _T_91 & _T_100; 
  assign _T_102 = _T_98 & _T_101; 
  assign _T_103 = _T_94 | _T_102; 
  assign _T_104 = _T_91 & _T_99; 
  assign _T_105 = _T_98 & _T_104; 
  assign _T_106 = _T_94 | _T_105; 
  assign _T_107 = _T_90 & _T_100; 
  assign _T_108 = _T_98 & _T_107; 
  assign _T_109 = _T_97 | _T_108; 
  assign _T_110 = _T_90 & _T_99; 
  assign _T_111 = _T_98 & _T_110; 
  assign _T_112 = _T_97 | _T_111; 
  assign _T_113 = _T_87[0]; 
  assign _T_114 = io_in_a_bits_address[0]; 
  assign _T_115 = _T_114 == 1'h0; 
  assign _T_116 = _T_101 & _T_115; 
  assign _T_117 = _T_113 & _T_116; 
  assign _T_118 = _T_103 | _T_117; 
  assign _T_119 = _T_101 & _T_114; 
  assign _T_120 = _T_113 & _T_119; 
  assign _T_121 = _T_103 | _T_120; 
  assign _T_122 = _T_104 & _T_115; 
  assign _T_123 = _T_113 & _T_122; 
  assign _T_124 = _T_106 | _T_123; 
  assign _T_125 = _T_104 & _T_114; 
  assign _T_126 = _T_113 & _T_125; 
  assign _T_127 = _T_106 | _T_126; 
  assign _T_128 = _T_107 & _T_115; 
  assign _T_129 = _T_113 & _T_128; 
  assign _T_130 = _T_109 | _T_129; 
  assign _T_131 = _T_107 & _T_114; 
  assign _T_132 = _T_113 & _T_131; 
  assign _T_133 = _T_109 | _T_132; 
  assign _T_134 = _T_110 & _T_115; 
  assign _T_135 = _T_113 & _T_134; 
  assign _T_136 = _T_112 | _T_135; 
  assign _T_137 = _T_110 & _T_114; 
  assign _T_138 = _T_113 & _T_137; 
  assign _T_139 = _T_112 | _T_138; 
  assign _T_146 = {_T_139,_T_136,_T_133,_T_130,_T_127,_T_124,_T_121,_T_118}; 
  assign _T_277 = io_in_a_bits_opcode == 3'h6; 
  assign _T_279 = io_in_a_bits_address ^ 32'h80000000; 
  assign _T_280 = {1'b0,$signed(_T_279)}; 
  assign _T_281 = $signed(_T_280) & $signed(-33'sh80000000); 
  assign _T_282 = $signed(_T_281); 
  assign _T_283 = $signed(_T_282) == $signed(33'sh0); 
  assign _T_288 = reset == 1'h0; 
  assign _T_355 = io_in_a_bits_size <= 3'h6; 
  assign _T_357 = _T_8 ? _T_355 : 1'h0; 
  assign _T_374 = _T_357 | reset; 
  assign _T_375 = _T_374 == 1'h0; 
  assign _T_377 = _T_76 | reset; 
  assign _T_378 = _T_377 == 1'h0; 
  assign _T_381 = _T_88 | reset; 
  assign _T_382 = _T_381 == 1'h0; 
  assign _T_384 = _T_82 | reset; 
  assign _T_385 = _T_384 == 1'h0; 
  assign _T_386 = io_in_a_bits_param <= 3'h2; 
  assign _T_388 = _T_386 | reset; 
  assign _T_389 = _T_388 == 1'h0; 
  assign _T_390 = ~ io_in_a_bits_mask; 
  assign _T_391 = _T_390 == 8'h0; 
  assign _T_393 = _T_391 | reset; 
  assign _T_394 = _T_393 == 1'h0; 
  assign _T_395 = io_in_a_bits_corrupt == 1'h0; 
  assign _T_397 = _T_395 | reset; 
  assign _T_398 = _T_397 == 1'h0; 
  assign _T_399 = io_in_a_bits_opcode == 3'h7; 
  assign _T_512 = io_in_a_bits_param != 3'h0; 
  assign _T_514 = _T_512 | reset; 
  assign _T_515 = _T_514 == 1'h0; 
  assign _T_525 = io_in_a_bits_opcode == 3'h4; 
  assign _T_535 = _T_355 & _T_283; 
  assign _T_538 = _T_535 | reset; 
  assign _T_539 = _T_538 == 1'h0; 
  assign _T_546 = io_in_a_bits_param == 3'h0; 
  assign _T_548 = _T_546 | reset; 
  assign _T_549 = _T_548 == 1'h0; 
  assign _T_550 = io_in_a_bits_mask == _T_146; 
  assign _T_552 = _T_550 | reset; 
  assign _T_553 = _T_552 == 1'h0; 
  assign _T_558 = io_in_a_bits_opcode == 3'h0; 
  assign _T_587 = io_in_a_bits_opcode == 3'h1; 
  assign _T_612 = ~ _T_146; 
  assign _T_613 = io_in_a_bits_mask & _T_612; 
  assign _T_614 = _T_613 == 8'h0; 
  assign _T_616 = _T_614 | reset; 
  assign _T_617 = _T_616 == 1'h0; 
  assign _T_618 = io_in_a_bits_opcode == 3'h2; 
  assign _T_636 = io_in_a_bits_param <= 3'h4; 
  assign _T_638 = _T_636 | reset; 
  assign _T_639 = _T_638 == 1'h0; 
  assign _T_644 = io_in_a_bits_opcode == 3'h3; 
  assign _T_662 = io_in_a_bits_param <= 3'h3; 
  assign _T_664 = _T_662 | reset; 
  assign _T_665 = _T_664 == 1'h0; 
  assign _T_670 = io_in_a_bits_opcode == 3'h5; 
  assign _T_696 = io_in_d_bits_opcode <= 3'h6; 
  assign _T_698 = _T_696 | reset; 
  assign _T_699 = _T_698 == 1'h0; 
  assign _T_702 = io_in_d_bits_source[6:4]; 
  assign _T_703 = _T_702 == 3'h0; 
  assign _T_711 = _T_702 == 3'h1; 
  assign _T_719 = _T_702 == 3'h2; 
  assign _T_727 = _T_702 == 3'h3; 
  assign _T_735 = _T_702 == 3'h4; 
  assign _T_743 = _T_702 == 3'h5; 
  assign _T_751 = _T_702 == 3'h6; 
  assign _T_759 = _T_702 == 3'h7; 
  assign _T_765 = _T_703 | _T_711; 
  assign _T_766 = _T_765 | _T_719; 
  assign _T_767 = _T_766 | _T_727; 
  assign _T_768 = _T_767 | _T_735; 
  assign _T_769 = _T_768 | _T_743; 
  assign _T_770 = _T_769 | _T_751; 
  assign _T_771 = _T_770 | _T_759; 
  assign _T_773 = io_in_d_bits_opcode == 3'h6; 
  assign _T_775 = _T_771 | reset; 
  assign _T_776 = _T_775 == 1'h0; 
  assign _T_777 = io_in_d_bits_size >= 3'h3; 
  assign _T_779 = _T_777 | reset; 
  assign _T_780 = _T_779 == 1'h0; 
  assign _T_785 = io_in_d_bits_corrupt == 1'h0; 
  assign _T_787 = _T_785 | reset; 
  assign _T_788 = _T_787 == 1'h0; 
  assign _T_789 = io_in_d_bits_denied == 1'h0; 
  assign _T_791 = _T_789 | reset; 
  assign _T_792 = _T_791 == 1'h0; 
  assign _T_793 = io_in_d_bits_opcode == 3'h4; 
  assign _T_821 = io_in_d_bits_opcode == 3'h5; 
  assign _T_841 = _T_789 | io_in_d_bits_corrupt; 
  assign _T_843 = _T_841 | reset; 
  assign _T_844 = _T_843 == 1'h0; 
  assign _T_850 = io_in_d_bits_opcode == 3'h0; 
  assign _T_867 = io_in_d_bits_opcode == 3'h1; 
  assign _T_885 = io_in_d_bits_opcode == 3'h2; 
  assign _T_914 = io_in_a_ready & io_in_a_valid; 
  assign _T_919 = _T_80[5:3]; 
  assign _T_920 = io_in_a_bits_opcode[2]; 
  assign _T_921 = _T_920 == 1'h0; 
  assign _T_925 = _T_923 - 3'h1; 
  assign _T_926 = _T_923 == 3'h0; 
  assign _T_939 = _T_926 == 1'h0; 
  assign _T_940 = io_in_a_valid & _T_939; 
  assign _T_941 = io_in_a_bits_opcode == _T_934; 
  assign _T_943 = _T_941 | reset; 
  assign _T_944 = _T_943 == 1'h0; 
  assign _T_945 = io_in_a_bits_param == _T_935; 
  assign _T_947 = _T_945 | reset; 
  assign _T_948 = _T_947 == 1'h0; 
  assign _T_949 = io_in_a_bits_size == _T_936; 
  assign _T_951 = _T_949 | reset; 
  assign _T_952 = _T_951 == 1'h0; 
  assign _T_953 = io_in_a_bits_source == _T_937; 
  assign _T_955 = _T_953 | reset; 
  assign _T_956 = _T_955 == 1'h0; 
  assign _T_957 = io_in_a_bits_address == _T_938; 
  assign _T_959 = _T_957 | reset; 
  assign _T_960 = _T_959 == 1'h0; 
  assign _T_962 = _T_914 & _T_926; 
  assign _T_963 = io_in_d_ready & io_in_d_valid; 
  assign _T_965 = 13'h3f << io_in_d_bits_size; 
  assign _T_966 = _T_965[5:0]; 
  assign _T_967 = ~ _T_966; 
  assign _T_968 = _T_967[5:3]; 
  assign _T_969 = io_in_d_bits_opcode[0]; 
  assign _T_973 = _T_971 - 3'h1; 
  assign _T_974 = _T_971 == 3'h0; 
  assign _T_988 = _T_974 == 1'h0; 
  assign _T_989 = io_in_d_valid & _T_988; 
  assign _T_990 = io_in_d_bits_opcode == _T_982; 
  assign _T_992 = _T_990 | reset; 
  assign _T_993 = _T_992 == 1'h0; 
  assign _T_998 = io_in_d_bits_size == _T_984; 
  assign _T_1000 = _T_998 | reset; 
  assign _T_1001 = _T_1000 == 1'h0; 
  assign _T_1002 = io_in_d_bits_source == _T_985; 
  assign _T_1004 = _T_1002 | reset; 
  assign _T_1005 = _T_1004 == 1'h0; 
  assign _T_1010 = io_in_d_bits_denied == _T_987; 
  assign _T_1012 = _T_1010 | reset; 
  assign _T_1013 = _T_1012 == 1'h0; 
  assign _T_1015 = _T_963 & _T_974; 
  assign _T_1028 = _T_1026 - 3'h1; 
  assign _T_1029 = _T_1026 == 3'h0; 
  assign _T_1047 = _T_1045 - 3'h1; 
  assign _T_1048 = _T_1045 == 3'h0; 
  assign _T_1058 = _T_914 & _T_1029; 
  assign _T_1060 = 128'h1 << io_in_a_bits_source; 
  assign _T_1061 = _T_1016 >> io_in_a_bits_source; 
  assign _T_1062 = _T_1061[0]; 
  assign _T_1063 = _T_1062 == 1'h0; 
  assign _T_1065 = _T_1063 | reset; 
  assign _T_1066 = _T_1065 == 1'h0; 
  assign _GEN_15 = _T_1058 ? _T_1060 : 128'h0; 
  assign _T_1070 = _T_963 & _T_1048; 
  assign _T_1072 = _T_773 == 1'h0; 
  assign _T_1073 = _T_1070 & _T_1072; 
  assign _T_1074 = 128'h1 << io_in_d_bits_source; 
  assign _T_1075 = _GEN_15 | _T_1016; 
  assign _T_1076 = _T_1075 >> io_in_d_bits_source; 
  assign _T_1077 = _T_1076[0]; 
  assign _T_1079 = _T_1077 | reset; 
  assign _T_1080 = _T_1079 == 1'h0; 
  assign _GEN_16 = _T_1073 ? _T_1074 : 128'h0; 
  assign _T_1081 = _GEN_15 != _GEN_16; 
  assign _T_1082 = _GEN_15 != 128'h0; 
  assign _T_1083 = _T_1082 == 1'h0; 
  assign _T_1084 = _T_1081 | _T_1083; 
  assign _T_1086 = _T_1084 | reset; 
  assign _T_1087 = _T_1086 == 1'h0; 
  assign _T_1088 = _T_1016 | _GEN_15; 
  assign _T_1089 = ~ _GEN_16; 
  assign _T_1090 = _T_1088 & _T_1089; 
  assign _T_1092 = _T_1016 != 128'h0; 
  assign _T_1093 = _T_1092 == 1'h0; 
  assign _T_1094 = plusarg_reader_out == 32'h0; 
  assign _T_1095 = _T_1093 | _T_1094; 
  assign _T_1096 = _T_1091 < plusarg_reader_out; 
  assign _T_1097 = _T_1095 | _T_1096; 
  assign _T_1099 = _T_1097 | reset; 
  assign _T_1100 = _T_1099 == 1'h0; 
  assign _T_1102 = _T_1091 + 32'h1; 
  assign _T_1105 = _T_914 | _T_963; 
  assign _GEN_19 = io_in_a_valid & _T_277; 
  assign _GEN_35 = io_in_a_valid & _T_399; 
  assign _GEN_53 = io_in_a_valid & _T_525; 
  assign _GEN_65 = io_in_a_valid & _T_558; 
  assign _GEN_75 = io_in_a_valid & _T_587; 
  assign _GEN_85 = io_in_a_valid & _T_618; 
  assign _GEN_95 = io_in_a_valid & _T_644; 
  assign _GEN_105 = io_in_a_valid & _T_670; 
  assign _GEN_115 = io_in_d_valid & _T_773; 
  assign _GEN_123 = io_in_d_valid & _T_793; 
  assign _GEN_131 = io_in_d_valid & _T_821; 
  assign _GEN_139 = io_in_d_valid & _T_850; 
  assign _GEN_143 = io_in_d_valid & _T_867; 
  assign _GEN_147 = io_in_d_valid & _T_885; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_923 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_934 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_935 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_936 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_937 = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_938 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_971 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_982 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_984 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_985 = _RAND_9[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_987 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {4{`RANDOM}};
  _T_1016 = _RAND_11[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_1026 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_1045 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_1091 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_923 <= 3'h0;
    end else begin
      if (_T_914) begin
        if (_T_926) begin
          if (_T_921) begin
            _T_923 <= _T_919;
          end else begin
            _T_923 <= 3'h0;
          end
        end else begin
          _T_923 <= _T_925;
        end
      end
    end
    if (_T_962) begin
      _T_934 <= io_in_a_bits_opcode;
    end
    if (_T_962) begin
      _T_935 <= io_in_a_bits_param;
    end
    if (_T_962) begin
      _T_936 <= io_in_a_bits_size;
    end
    if (_T_962) begin
      _T_937 <= io_in_a_bits_source;
    end
    if (_T_962) begin
      _T_938 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_971 <= 3'h0;
    end else begin
      if (_T_963) begin
        if (_T_974) begin
          if (_T_969) begin
            _T_971 <= _T_968;
          end else begin
            _T_971 <= 3'h0;
          end
        end else begin
          _T_971 <= _T_973;
        end
      end
    end
    if (_T_1015) begin
      _T_982 <= io_in_d_bits_opcode;
    end
    if (_T_1015) begin
      _T_984 <= io_in_d_bits_size;
    end
    if (_T_1015) begin
      _T_985 <= io_in_d_bits_source;
    end
    if (_T_1015) begin
      _T_987 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_1016 <= 128'h0;
    end else begin
      _T_1016 <= _T_1090;
    end
    if (reset) begin
      _T_1026 <= 3'h0;
    end else begin
      if (_T_914) begin
        if (_T_1029) begin
          if (_T_921) begin
            _T_1026 <= _T_919;
          end else begin
            _T_1026 <= 3'h0;
          end
        end else begin
          _T_1026 <= _T_1028;
        end
      end
    end
    if (reset) begin
      _T_1045 <= 3'h0;
    end else begin
      if (_T_963) begin
        if (_T_1048) begin
          if (_T_969) begin
            _T_1045 <= _T_968;
          end else begin
            _T_1045 <= 3'h0;
          end
        end else begin
          _T_1045 <= _T_1047;
        end
      end
    end
    if (reset) begin
      _T_1091 <= 32'h0;
    end else begin
      if (_T_1105) begin
        _T_1091 <= 32'h0;
      end else begin
        _T_1091 <= _T_1102;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel has invalid opcode (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:39 assert (TLMessages.isA(bundle.opcode), \"'A' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:46 assert (visible(edge.address(bundle), bundle.source, edge), \"'A' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_288) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_288) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_375) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_375) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_378) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_378) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_382) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_382) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_385) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_389) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_389) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_394) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_394) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_398) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:56 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_398) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_288) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_288) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_375) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_375) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_378) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_378) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_382) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_382) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_385) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_389) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_389) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_515) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_515) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_394) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_394) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_398) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:68 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_398) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_539) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_539) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_378) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_378) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_385) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_549) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_549) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_553) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_553) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_398) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:77 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_53 & _T_398) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_539) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_539) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_378) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_378) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_385) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_549) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_549) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_65 & _T_553) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_65 & _T_553) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_539) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_539) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_378) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_378) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_385) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_549) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_549) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_617) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_617) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_288) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_288) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_378) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_378) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_385) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_639) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_639) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_553) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_85 & _T_553) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_288) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_288) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_378) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_378) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_385) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_665) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_665) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_95 & _T_553) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_95 & _T_553) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_288) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_288) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_378) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_378) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_385) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_385) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_553) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_553) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_398) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:117 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_398) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_699) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_699) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_776) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_776) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_780) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_780) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_788) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_788) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_115 & _T_792) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_115 & _T_792) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_776) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_776) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_288) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:285 assert (sink_ok, \"'D' channel Grant carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_288) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_780) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_780) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_788) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_123 & _T_788) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is denied (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:290 assert (deny_put_ok || !bundle.denied, \"'D' channel Grant is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_776) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_776) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_288) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:295 assert (sink_ok, \"'D' channel GrantData carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_288) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_780) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_780) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_844) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_844) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:300 assert (deny_get_ok || !bundle.denied, \"'D' channel GrantData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_139 & _T_776) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_139 & _T_776) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_139 & _T_788) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_139 & _T_788) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is denied (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:308 assert (deny_put_ok || !bundle.denied, \"'D' channel AccessAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & _T_776) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & _T_776) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & _T_844) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & _T_844) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:316 assert (deny_get_ok || !bundle.denied, \"'D' channel AccessAckData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_147 & _T_776) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_147 & _T_776) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_147 & _T_788) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_147 & _T_788) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is denied (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:324 assert (deny_put_ok || !bundle.denied, \"'D' channel HintAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel valid and not TL-C (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:341 assert (!bundle.b.valid, \"'B' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel valid and not TL-C (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:342 assert (!bundle.c.valid, \"'C' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel valid and not TL-C (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:343 assert (!bundle.e.valid, \"'E' channel valid and not TL-C\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_940 & _T_944) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_940 & _T_944) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_940 & _T_948) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_940 & _T_948) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_940 & _T_952) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_940 & _T_952) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_940 & _T_956) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_940 & _T_956) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_940 & _T_960) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_940 & _T_960) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_989 & _T_993) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_989 & _T_993) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_989 & _T_1001) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_989 & _T_1001) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_989 & _T_1005) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_989 & _T_1005) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_989 & _T_1013) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_989 & _T_1013) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1058 & _T_1066) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1058 & _T_1066) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1073 & _T_1080) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1073 & _T_1080) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1087) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1087) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1100) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at ChiplinkTest.scala:178:90)\n    at Monitor.scala:479 assert (!inflight.orR || limit === UInt(0) || watchdog < limit, \"TileLink timeout expired\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1100) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLMonitor( 
  input         clock, 
  input         reset, 
  input         io_in_a_ready, 
  input         io_in_a_valid, 
  input  [2:0]  io_in_a_bits_opcode, 
  input  [2:0]  io_in_a_bits_param, 
  input  [3:0]  io_in_a_bits_size, 
  input  [6:0]  io_in_a_bits_source, 
  input  [31:0] io_in_a_bits_address, 
  input  [7:0]  io_in_a_bits_mask, 
  input         io_in_a_bits_corrupt, 
  input         io_in_c_ready, 
  input         io_in_c_valid, 
  input  [2:0]  io_in_c_bits_opcode, 
  input  [2:0]  io_in_c_bits_param, 
  input  [3:0]  io_in_c_bits_size, 
  input  [6:0]  io_in_c_bits_source, 
  input  [31:0] io_in_c_bits_address, 
  input         io_in_c_bits_corrupt, 
  input         io_in_d_ready, 
  input         io_in_d_valid, 
  input  [2:0]  io_in_d_bits_opcode, 
  input  [1:0]  io_in_d_bits_param, 
  input  [3:0]  io_in_d_bits_size, 
  input  [6:0]  io_in_d_bits_source, 
  input         io_in_d_bits_sink, 
  input         io_in_d_bits_denied, 
  input         io_in_d_bits_corrupt, 
  input         io_in_e_ready, 
  input         io_in_e_valid, 
  input         io_in_e_bits_sink 
);
  wire [31:0] plusarg_reader_out; 
  wire [2:0] _T_7; 
  wire  _T_8; 
  wire  _T_16; 
  wire  _T_24; 
  wire  _T_32; 
  wire  _T_40; 
  wire  _T_48; 
  wire  _T_56; 
  wire  _T_64; 
  wire  _T_70; 
  wire  _T_71; 
  wire  _T_72; 
  wire  _T_73; 
  wire  _T_74; 
  wire  _T_75; 
  wire  _T_76; 
  wire [22:0] _T_78; 
  wire [7:0] _T_79; 
  wire [7:0] _T_80; 
  wire [31:0] _GEN_33; 
  wire [31:0] _T_81; 
  wire  _T_82; 
  wire [1:0] _T_84; 
  wire [3:0] _T_85; 
  wire [2:0] _T_86; 
  wire [2:0] _T_87; 
  wire  _T_88; 
  wire  _T_89; 
  wire  _T_90; 
  wire  _T_91; 
  wire  _T_93; 
  wire  _T_94; 
  wire  _T_96; 
  wire  _T_97; 
  wire  _T_98; 
  wire  _T_99; 
  wire  _T_100; 
  wire  _T_101; 
  wire  _T_102; 
  wire  _T_103; 
  wire  _T_104; 
  wire  _T_105; 
  wire  _T_106; 
  wire  _T_107; 
  wire  _T_108; 
  wire  _T_109; 
  wire  _T_110; 
  wire  _T_111; 
  wire  _T_112; 
  wire  _T_113; 
  wire  _T_114; 
  wire  _T_115; 
  wire  _T_116; 
  wire  _T_117; 
  wire  _T_118; 
  wire  _T_119; 
  wire  _T_120; 
  wire  _T_121; 
  wire  _T_122; 
  wire  _T_123; 
  wire  _T_124; 
  wire  _T_125; 
  wire  _T_126; 
  wire  _T_127; 
  wire  _T_128; 
  wire  _T_129; 
  wire  _T_130; 
  wire  _T_131; 
  wire  _T_132; 
  wire  _T_133; 
  wire  _T_134; 
  wire  _T_135; 
  wire  _T_136; 
  wire  _T_137; 
  wire  _T_138; 
  wire  _T_139; 
  wire [7:0] _T_146; 
  wire  _T_277; 
  wire [31:0] _T_279; 
  wire [32:0] _T_280; 
  wire [32:0] _T_281; 
  wire [32:0] _T_282; 
  wire  _T_283; 
  wire [31:0] _T_284; 
  wire [32:0] _T_285; 
  wire [32:0] _T_286; 
  wire [32:0] _T_287; 
  wire  _T_288; 
  wire  _T_289; 
  wire  _T_292; 
  wire [31:0] _T_295; 
  wire [32:0] _T_296; 
  wire [32:0] _T_297; 
  wire [32:0] _T_298; 
  wire  _T_299; 
  wire  _T_300; 
  wire  _T_304; 
  wire  _T_305; 
  wire  _T_374; 
  wire  _T_391; 
  wire  _T_392; 
  wire  _T_394; 
  wire  _T_395; 
  wire  _T_398; 
  wire  _T_399; 
  wire  _T_401; 
  wire  _T_402; 
  wire  _T_403; 
  wire  _T_405; 
  wire  _T_406; 
  wire [7:0] _T_407; 
  wire  _T_408; 
  wire  _T_410; 
  wire  _T_411; 
  wire  _T_412; 
  wire  _T_414; 
  wire  _T_415; 
  wire  _T_416; 
  wire  _T_546; 
  wire  _T_548; 
  wire  _T_549; 
  wire  _T_559; 
  wire  _T_580; 
  wire  _T_581; 
  wire  _T_584; 
  wire  _T_585; 
  wire  _T_592; 
  wire  _T_594; 
  wire  _T_595; 
  wire  _T_596; 
  wire  _T_598; 
  wire  _T_599; 
  wire  _T_604; 
  wire  _T_619; 
  wire  _T_620; 
  wire  _T_622; 
  wire  _T_630; 
  wire  _T_632; 
  wire  _T_634; 
  wire  _T_635; 
  wire  _T_650; 
  wire [7:0] _T_692; 
  wire [7:0] _T_693; 
  wire  _T_694; 
  wire  _T_696; 
  wire  _T_697; 
  wire  _T_698; 
  wire  _T_733; 
  wire  _T_735; 
  wire  _T_736; 
  wire  _T_741; 
  wire  _T_776; 
  wire  _T_778; 
  wire  _T_779; 
  wire  _T_784; 
  wire  _T_827; 
  wire  _T_829; 
  wire  _T_830; 
  wire [2:0] _T_833; 
  wire  _T_834; 
  wire  _T_842; 
  wire  _T_850; 
  wire  _T_858; 
  wire  _T_866; 
  wire  _T_874; 
  wire  _T_882; 
  wire  _T_890; 
  wire  _T_896; 
  wire  _T_897; 
  wire  _T_898; 
  wire  _T_899; 
  wire  _T_900; 
  wire  _T_901; 
  wire  _T_902; 
  wire  _T_903; 
  wire  _T_904; 
  wire  _T_906; 
  wire  _T_907; 
  wire  _T_908; 
  wire  _T_910; 
  wire  _T_911; 
  wire  _T_912; 
  wire  _T_914; 
  wire  _T_915; 
  wire  _T_916; 
  wire  _T_918; 
  wire  _T_919; 
  wire  _T_920; 
  wire  _T_922; 
  wire  _T_923; 
  wire  _T_924; 
  wire  _T_929; 
  wire  _T_930; 
  wire  _T_935; 
  wire  _T_937; 
  wire  _T_938; 
  wire  _T_939; 
  wire  _T_941; 
  wire  _T_942; 
  wire  _T_952; 
  wire  _T_972; 
  wire  _T_974; 
  wire  _T_975; 
  wire  _T_981; 
  wire  _T_998; 
  wire  _T_1016; 
  wire [2:0] _T_1584; 
  wire  _T_1585; 
  wire  _T_1593; 
  wire  _T_1601; 
  wire  _T_1609; 
  wire  _T_1617; 
  wire  _T_1625; 
  wire  _T_1633; 
  wire  _T_1641; 
  wire  _T_1647; 
  wire  _T_1648; 
  wire  _T_1649; 
  wire  _T_1650; 
  wire  _T_1651; 
  wire  _T_1652; 
  wire  _T_1653; 
  wire [22:0] _T_1655; 
  wire [7:0] _T_1656; 
  wire [7:0] _T_1657; 
  wire [31:0] _GEN_34; 
  wire [31:0] _T_1658; 
  wire  _T_1659; 
  wire [31:0] _T_1660; 
  wire [32:0] _T_1661; 
  wire [32:0] _T_1662; 
  wire [32:0] _T_1663; 
  wire  _T_1664; 
  wire [31:0] _T_1665; 
  wire [32:0] _T_1666; 
  wire [32:0] _T_1667; 
  wire [32:0] _T_1668; 
  wire  _T_1669; 
  wire [31:0] _T_1670; 
  wire [32:0] _T_1671; 
  wire [32:0] _T_1672; 
  wire [32:0] _T_1673; 
  wire  _T_1674; 
  wire  _T_1676; 
  wire  _T_1677; 
  wire  _T_1808; 
  wire  _T_1810; 
  wire  _T_1811; 
  wire  _T_1813; 
  wire  _T_1814; 
  wire  _T_1815; 
  wire  _T_1817; 
  wire  _T_1818; 
  wire  _T_1820; 
  wire  _T_1821; 
  wire  _T_1822; 
  wire  _T_1824; 
  wire  _T_1825; 
  wire  _T_1826; 
  wire  _T_1828; 
  wire  _T_1829; 
  wire  _T_1830; 
  wire  _T_1848; 
  wire  _T_1863; 
  wire  _T_1871; 
  wire  _T_1875; 
  wire  _T_1876; 
  wire  _T_1945; 
  wire  _T_1962; 
  wire  _T_1963; 
  wire  _T_1974; 
  wire  _T_1976; 
  wire  _T_1977; 
  wire  _T_1982; 
  wire  _T_2112; 
  wire  _T_2122; 
  wire  _T_2124; 
  wire  _T_2125; 
  wire  _T_2130; 
  wire  _T_2144; 
  wire  _T_2162; 
  wire  _T_2164; 
  wire  _T_2165; 
  wire  _T_2166; 
  wire [4:0] _T_2171; 
  wire  _T_2172; 
  wire  _T_2173; 
  reg [4:0] _T_2175; 
  reg [31:0] _RAND_0;
  wire [4:0] _T_2177; 
  wire  _T_2178; 
  reg [2:0] _T_2186; 
  reg [31:0] _RAND_1;
  reg [2:0] _T_2187; 
  reg [31:0] _RAND_2;
  reg [3:0] _T_2188; 
  reg [31:0] _RAND_3;
  reg [6:0] _T_2189; 
  reg [31:0] _RAND_4;
  reg [31:0] _T_2190; 
  reg [31:0] _RAND_5;
  wire  _T_2191; 
  wire  _T_2192; 
  wire  _T_2193; 
  wire  _T_2195; 
  wire  _T_2196; 
  wire  _T_2197; 
  wire  _T_2199; 
  wire  _T_2200; 
  wire  _T_2201; 
  wire  _T_2203; 
  wire  _T_2204; 
  wire  _T_2205; 
  wire  _T_2207; 
  wire  _T_2208; 
  wire  _T_2209; 
  wire  _T_2211; 
  wire  _T_2212; 
  wire  _T_2214; 
  wire  _T_2215; 
  wire [22:0] _T_2217; 
  wire [7:0] _T_2218; 
  wire [7:0] _T_2219; 
  wire [4:0] _T_2220; 
  wire  _T_2221; 
  reg [4:0] _T_2223; 
  reg [31:0] _RAND_6;
  wire [4:0] _T_2225; 
  wire  _T_2226; 
  reg [2:0] _T_2234; 
  reg [31:0] _RAND_7;
  reg [1:0] _T_2235; 
  reg [31:0] _RAND_8;
  reg [3:0] _T_2236; 
  reg [31:0] _RAND_9;
  reg [6:0] _T_2237; 
  reg [31:0] _RAND_10;
  reg  _T_2238; 
  reg [31:0] _RAND_11;
  reg  _T_2239; 
  reg [31:0] _RAND_12;
  wire  _T_2240; 
  wire  _T_2241; 
  wire  _T_2242; 
  wire  _T_2244; 
  wire  _T_2245; 
  wire  _T_2246; 
  wire  _T_2248; 
  wire  _T_2249; 
  wire  _T_2250; 
  wire  _T_2252; 
  wire  _T_2253; 
  wire  _T_2254; 
  wire  _T_2256; 
  wire  _T_2257; 
  wire  _T_2258; 
  wire  _T_2260; 
  wire  _T_2261; 
  wire  _T_2262; 
  wire  _T_2264; 
  wire  _T_2265; 
  wire  _T_2267; 
  wire  _T_2317; 
  wire [4:0] _T_2322; 
  wire  _T_2323; 
  reg [4:0] _T_2325; 
  reg [31:0] _RAND_13;
  wire [4:0] _T_2327; 
  wire  _T_2328; 
  reg [2:0] _T_2336; 
  reg [31:0] _RAND_14;
  reg [2:0] _T_2337; 
  reg [31:0] _RAND_15;
  reg [3:0] _T_2338; 
  reg [31:0] _RAND_16;
  reg [6:0] _T_2339; 
  reg [31:0] _RAND_17;
  reg [31:0] _T_2340; 
  reg [31:0] _RAND_18;
  wire  _T_2341; 
  wire  _T_2342; 
  wire  _T_2343; 
  wire  _T_2345; 
  wire  _T_2346; 
  wire  _T_2347; 
  wire  _T_2349; 
  wire  _T_2350; 
  wire  _T_2351; 
  wire  _T_2353; 
  wire  _T_2354; 
  wire  _T_2355; 
  wire  _T_2357; 
  wire  _T_2358; 
  wire  _T_2359; 
  wire  _T_2361; 
  wire  _T_2362; 
  wire  _T_2364; 
  reg [127:0] _T_2365; 
  reg [127:0] _RAND_19;
  reg [4:0] _T_2375; 
  reg [31:0] _RAND_20;
  wire [4:0] _T_2377; 
  wire  _T_2378; 
  reg [4:0] _T_2394; 
  reg [31:0] _RAND_21;
  wire [4:0] _T_2396; 
  wire  _T_2397; 
  wire  _T_2407; 
  wire [127:0] _T_2409; 
  wire [127:0] _T_2410; 
  wire  _T_2411; 
  wire  _T_2412; 
  wire  _T_2414; 
  wire  _T_2415; 
  wire [127:0] _GEN_27; 
  wire  _T_2419; 
  wire  _T_2421; 
  wire  _T_2422; 
  wire [127:0] _T_2423; 
  wire [127:0] _T_2424; 
  wire [127:0] _T_2425; 
  wire  _T_2426; 
  wire  _T_2428; 
  wire  _T_2429; 
  wire [127:0] _GEN_28; 
  wire  _T_2430; 
  wire  _T_2431; 
  wire  _T_2432; 
  wire  _T_2433; 
  wire  _T_2435; 
  wire  _T_2436; 
  wire [127:0] _T_2437; 
  wire [127:0] _T_2438; 
  wire [127:0] _T_2439; 
  reg [31:0] _T_2440; 
  reg [31:0] _RAND_22;
  wire  _T_2441; 
  wire  _T_2442; 
  wire  _T_2443; 
  wire  _T_2444; 
  wire  _T_2445; 
  wire  _T_2446; 
  wire  _T_2448; 
  wire  _T_2449; 
  wire [31:0] _T_2451; 
  wire  _T_2454; 
  reg  _T_2455; 
  reg [31:0] _RAND_23;
  reg [4:0] _T_2464; 
  reg [31:0] _RAND_24;
  wire [4:0] _T_2466; 
  wire  _T_2467; 
  wire  _T_2477; 
  wire  _T_2478; 
  wire  _T_2479; 
  wire  _T_2480; 
  wire  _T_2481; 
  wire  _T_2482; 
  wire [1:0] _T_2483; 
  wire  _T_2484; 
  wire  _T_2486; 
  wire  _T_2488; 
  wire  _T_2489; 
  wire [1:0] _GEN_31; 
  wire  _T_2491; 
  wire [1:0] _T_2494; 
  wire  _T_2475; 
  wire  _T_2495; 
  wire  _T_2496; 
  wire  _T_2499; 
  wire  _T_2500; 
  wire [1:0] _GEN_32; 
  wire  _T_2501; 
  wire  _T_2490; 
  wire  _T_2502; 
  wire  _T_2503; 
  wire  _GEN_35; 
  wire  _GEN_51; 
  wire  _GEN_69; 
  wire  _GEN_81; 
  wire  _GEN_91; 
  wire  _GEN_101; 
  wire  _GEN_111; 
  wire  _GEN_121; 
  wire  _GEN_131; 
  wire  _GEN_141; 
  wire  _GEN_153; 
  wire  _GEN_165; 
  wire  _GEN_171; 
  wire  _GEN_177; 
  wire  _GEN_183; 
  wire  _GEN_195; 
  wire  _GEN_205; 
  wire  _GEN_219; 
  wire  _GEN_231; 
  wire  _GEN_241; 
  wire  _GEN_249; 
  dual_plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0)) plusarg_reader ( 
    .out(plusarg_reader_out)
  );
  assign _T_7 = io_in_a_bits_source[6:4]; 
  assign _T_8 = _T_7 == 3'h0; 
  assign _T_16 = _T_7 == 3'h1; 
  assign _T_24 = _T_7 == 3'h2; 
  assign _T_32 = _T_7 == 3'h3; 
  assign _T_40 = _T_7 == 3'h4; 
  assign _T_48 = _T_7 == 3'h5; 
  assign _T_56 = _T_7 == 3'h6; 
  assign _T_64 = _T_7 == 3'h7; 
  assign _T_70 = _T_8 | _T_16; 
  assign _T_71 = _T_70 | _T_24; 
  assign _T_72 = _T_71 | _T_32; 
  assign _T_73 = _T_72 | _T_40; 
  assign _T_74 = _T_73 | _T_48; 
  assign _T_75 = _T_74 | _T_56; 
  assign _T_76 = _T_75 | _T_64; 
  assign _T_78 = 23'hff << io_in_a_bits_size; 
  assign _T_79 = _T_78[7:0]; 
  assign _T_80 = ~ _T_79; 
  assign _GEN_33 = {{24'd0}, _T_80}; 
  assign _T_81 = io_in_a_bits_address & _GEN_33; 
  assign _T_82 = _T_81 == 32'h0; 
  assign _T_84 = io_in_a_bits_size[1:0]; 
  assign _T_85 = 4'h1 << _T_84; 
  assign _T_86 = _T_85[2:0]; 
  assign _T_87 = _T_86 | 3'h1; 
  assign _T_88 = io_in_a_bits_size >= 4'h3; 
  assign _T_89 = _T_87[2]; 
  assign _T_90 = io_in_a_bits_address[2]; 
  assign _T_91 = _T_90 == 1'h0; 
  assign _T_93 = _T_89 & _T_91; 
  assign _T_94 = _T_88 | _T_93; 
  assign _T_96 = _T_89 & _T_90; 
  assign _T_97 = _T_88 | _T_96; 
  assign _T_98 = _T_87[1]; 
  assign _T_99 = io_in_a_bits_address[1]; 
  assign _T_100 = _T_99 == 1'h0; 
  assign _T_101 = _T_91 & _T_100; 
  assign _T_102 = _T_98 & _T_101; 
  assign _T_103 = _T_94 | _T_102; 
  assign _T_104 = _T_91 & _T_99; 
  assign _T_105 = _T_98 & _T_104; 
  assign _T_106 = _T_94 | _T_105; 
  assign _T_107 = _T_90 & _T_100; 
  assign _T_108 = _T_98 & _T_107; 
  assign _T_109 = _T_97 | _T_108; 
  assign _T_110 = _T_90 & _T_99; 
  assign _T_111 = _T_98 & _T_110; 
  assign _T_112 = _T_97 | _T_111; 
  assign _T_113 = _T_87[0]; 
  assign _T_114 = io_in_a_bits_address[0]; 
  assign _T_115 = _T_114 == 1'h0; 
  assign _T_116 = _T_101 & _T_115; 
  assign _T_117 = _T_113 & _T_116; 
  assign _T_118 = _T_103 | _T_117; 
  assign _T_119 = _T_101 & _T_114; 
  assign _T_120 = _T_113 & _T_119; 
  assign _T_121 = _T_103 | _T_120; 
  assign _T_122 = _T_104 & _T_115; 
  assign _T_123 = _T_113 & _T_122; 
  assign _T_124 = _T_106 | _T_123; 
  assign _T_125 = _T_104 & _T_114; 
  assign _T_126 = _T_113 & _T_125; 
  assign _T_127 = _T_106 | _T_126; 
  assign _T_128 = _T_107 & _T_115; 
  assign _T_129 = _T_113 & _T_128; 
  assign _T_130 = _T_109 | _T_129; 
  assign _T_131 = _T_107 & _T_114; 
  assign _T_132 = _T_113 & _T_131; 
  assign _T_133 = _T_109 | _T_132; 
  assign _T_134 = _T_110 & _T_115; 
  assign _T_135 = _T_113 & _T_134; 
  assign _T_136 = _T_112 | _T_135; 
  assign _T_137 = _T_110 & _T_114; 
  assign _T_138 = _T_113 & _T_137; 
  assign _T_139 = _T_112 | _T_138; 
  assign _T_146 = {_T_139,_T_136,_T_133,_T_130,_T_127,_T_124,_T_121,_T_118}; 
  assign _T_277 = io_in_a_bits_opcode == 3'h6; 
  assign _T_279 = io_in_a_bits_address ^ 32'h80000000; 
  assign _T_280 = {1'b0,$signed(_T_279)}; 
  assign _T_281 = $signed(_T_280) & $signed(-33'sh80000000); 
  assign _T_282 = $signed(_T_281); 
  assign _T_283 = $signed(_T_282) == $signed(33'sh0); 
  assign _T_284 = io_in_a_bits_address ^ 32'h40000000; 
  assign _T_285 = {1'b0,$signed(_T_284)}; 
  assign _T_286 = $signed(_T_285) & $signed(-33'sh20000000); 
  assign _T_287 = $signed(_T_286); 
  assign _T_288 = $signed(_T_287) == $signed(33'sh0); 
  assign _T_289 = _T_283 | _T_288; 
  assign _T_292 = io_in_a_bits_size <= 4'h6; 
  assign _T_295 = io_in_a_bits_address ^ 32'h10000000; 
  assign _T_296 = {1'b0,$signed(_T_295)}; 
  assign _T_297 = $signed(_T_296) & $signed(-33'sh10000000); 
  assign _T_298 = $signed(_T_297); 
  assign _T_299 = $signed(_T_298) == $signed(33'sh0); 
  assign _T_300 = _T_292 & _T_299; 
  assign _T_304 = _T_300 | reset; 
  assign _T_305 = _T_304 == 1'h0; 
  assign _T_374 = _T_8 ? _T_292 : 1'h0; 
  assign _T_391 = _T_374 | reset; 
  assign _T_392 = _T_391 == 1'h0; 
  assign _T_394 = _T_76 | reset; 
  assign _T_395 = _T_394 == 1'h0; 
  assign _T_398 = _T_88 | reset; 
  assign _T_399 = _T_398 == 1'h0; 
  assign _T_401 = _T_82 | reset; 
  assign _T_402 = _T_401 == 1'h0; 
  assign _T_403 = io_in_a_bits_param <= 3'h2; 
  assign _T_405 = _T_403 | reset; 
  assign _T_406 = _T_405 == 1'h0; 
  assign _T_407 = ~ io_in_a_bits_mask; 
  assign _T_408 = _T_407 == 8'h0; 
  assign _T_410 = _T_408 | reset; 
  assign _T_411 = _T_410 == 1'h0; 
  assign _T_412 = io_in_a_bits_corrupt == 1'h0; 
  assign _T_414 = _T_412 | reset; 
  assign _T_415 = _T_414 == 1'h0; 
  assign _T_416 = io_in_a_bits_opcode == 3'h7; 
  assign _T_546 = io_in_a_bits_param != 3'h0; 
  assign _T_548 = _T_546 | reset; 
  assign _T_549 = _T_548 == 1'h0; 
  assign _T_559 = io_in_a_bits_opcode == 3'h4; 
  assign _T_580 = _T_289 | _T_299; 
  assign _T_581 = _T_292 & _T_580; 
  assign _T_584 = _T_581 | reset; 
  assign _T_585 = _T_584 == 1'h0; 
  assign _T_592 = io_in_a_bits_param == 3'h0; 
  assign _T_594 = _T_592 | reset; 
  assign _T_595 = _T_594 == 1'h0; 
  assign _T_596 = io_in_a_bits_mask == _T_146; 
  assign _T_598 = _T_596 | reset; 
  assign _T_599 = _T_598 == 1'h0; 
  assign _T_604 = io_in_a_bits_opcode == 3'h0; 
  assign _T_619 = _T_283 | _T_299; 
  assign _T_620 = _T_292 & _T_619; 
  assign _T_622 = io_in_a_bits_size <= 4'h8; 
  assign _T_630 = _T_622 & _T_288; 
  assign _T_632 = _T_620 | _T_630; 
  assign _T_634 = _T_632 | reset; 
  assign _T_635 = _T_634 == 1'h0; 
  assign _T_650 = io_in_a_bits_opcode == 3'h1; 
  assign _T_692 = ~ _T_146; 
  assign _T_693 = io_in_a_bits_mask & _T_692; 
  assign _T_694 = _T_693 == 8'h0; 
  assign _T_696 = _T_694 | reset; 
  assign _T_697 = _T_696 == 1'h0; 
  assign _T_698 = io_in_a_bits_opcode == 3'h2; 
  assign _T_733 = io_in_a_bits_param <= 3'h4; 
  assign _T_735 = _T_733 | reset; 
  assign _T_736 = _T_735 == 1'h0; 
  assign _T_741 = io_in_a_bits_opcode == 3'h3; 
  assign _T_776 = io_in_a_bits_param <= 3'h3; 
  assign _T_778 = _T_776 | reset; 
  assign _T_779 = _T_778 == 1'h0; 
  assign _T_784 = io_in_a_bits_opcode == 3'h5; 
  assign _T_827 = io_in_d_bits_opcode <= 3'h6; 
  assign _T_829 = _T_827 | reset; 
  assign _T_830 = _T_829 == 1'h0; 
  assign _T_833 = io_in_d_bits_source[6:4]; 
  assign _T_834 = _T_833 == 3'h0; 
  assign _T_842 = _T_833 == 3'h1; 
  assign _T_850 = _T_833 == 3'h2; 
  assign _T_858 = _T_833 == 3'h3; 
  assign _T_866 = _T_833 == 3'h4; 
  assign _T_874 = _T_833 == 3'h5; 
  assign _T_882 = _T_833 == 3'h6; 
  assign _T_890 = _T_833 == 3'h7; 
  assign _T_896 = _T_834 | _T_842; 
  assign _T_897 = _T_896 | _T_850; 
  assign _T_898 = _T_897 | _T_858; 
  assign _T_899 = _T_898 | _T_866; 
  assign _T_900 = _T_899 | _T_874; 
  assign _T_901 = _T_900 | _T_882; 
  assign _T_902 = _T_901 | _T_890; 
  assign _T_903 = io_in_d_bits_sink < 1'h1; 
  assign _T_904 = io_in_d_bits_opcode == 3'h6; 
  assign _T_906 = _T_902 | reset; 
  assign _T_907 = _T_906 == 1'h0; 
  assign _T_908 = io_in_d_bits_size >= 4'h3; 
  assign _T_910 = _T_908 | reset; 
  assign _T_911 = _T_910 == 1'h0; 
  assign _T_912 = io_in_d_bits_param == 2'h0; 
  assign _T_914 = _T_912 | reset; 
  assign _T_915 = _T_914 == 1'h0; 
  assign _T_916 = io_in_d_bits_corrupt == 1'h0; 
  assign _T_918 = _T_916 | reset; 
  assign _T_919 = _T_918 == 1'h0; 
  assign _T_920 = io_in_d_bits_denied == 1'h0; 
  assign _T_922 = _T_920 | reset; 
  assign _T_923 = _T_922 == 1'h0; 
  assign _T_924 = io_in_d_bits_opcode == 3'h4; 
  assign _T_929 = _T_903 | reset; 
  assign _T_930 = _T_929 == 1'h0; 
  assign _T_935 = io_in_d_bits_param <= 2'h2; 
  assign _T_937 = _T_935 | reset; 
  assign _T_938 = _T_937 == 1'h0; 
  assign _T_939 = io_in_d_bits_param != 2'h2; 
  assign _T_941 = _T_939 | reset; 
  assign _T_942 = _T_941 == 1'h0; 
  assign _T_952 = io_in_d_bits_opcode == 3'h5; 
  assign _T_972 = _T_920 | io_in_d_bits_corrupt; 
  assign _T_974 = _T_972 | reset; 
  assign _T_975 = _T_974 == 1'h0; 
  assign _T_981 = io_in_d_bits_opcode == 3'h0; 
  assign _T_998 = io_in_d_bits_opcode == 3'h1; 
  assign _T_1016 = io_in_d_bits_opcode == 3'h2; 
  assign _T_1584 = io_in_c_bits_source[6:4]; 
  assign _T_1585 = _T_1584 == 3'h0; 
  assign _T_1593 = _T_1584 == 3'h1; 
  assign _T_1601 = _T_1584 == 3'h2; 
  assign _T_1609 = _T_1584 == 3'h3; 
  assign _T_1617 = _T_1584 == 3'h4; 
  assign _T_1625 = _T_1584 == 3'h5; 
  assign _T_1633 = _T_1584 == 3'h6; 
  assign _T_1641 = _T_1584 == 3'h7; 
  assign _T_1647 = _T_1585 | _T_1593; 
  assign _T_1648 = _T_1647 | _T_1601; 
  assign _T_1649 = _T_1648 | _T_1609; 
  assign _T_1650 = _T_1649 | _T_1617; 
  assign _T_1651 = _T_1650 | _T_1625; 
  assign _T_1652 = _T_1651 | _T_1633; 
  assign _T_1653 = _T_1652 | _T_1641; 
  assign _T_1655 = 23'hff << io_in_c_bits_size; 
  assign _T_1656 = _T_1655[7:0]; 
  assign _T_1657 = ~ _T_1656; 
  assign _GEN_34 = {{24'd0}, _T_1657}; 
  assign _T_1658 = io_in_c_bits_address & _GEN_34; 
  assign _T_1659 = _T_1658 == 32'h0; 
  assign _T_1660 = io_in_c_bits_address ^ 32'h80000000; 
  assign _T_1661 = {1'b0,$signed(_T_1660)}; 
  assign _T_1662 = $signed(_T_1661) & $signed(-33'sh80000000); 
  assign _T_1663 = $signed(_T_1662); 
  assign _T_1664 = $signed(_T_1663) == $signed(33'sh0); 
  assign _T_1665 = io_in_c_bits_address ^ 32'h40000000; 
  assign _T_1666 = {1'b0,$signed(_T_1665)}; 
  assign _T_1667 = $signed(_T_1666) & $signed(-33'sh20000000); 
  assign _T_1668 = $signed(_T_1667); 
  assign _T_1669 = $signed(_T_1668) == $signed(33'sh0); 
  assign _T_1670 = io_in_c_bits_address ^ 32'h10000000; 
  assign _T_1671 = {1'b0,$signed(_T_1670)}; 
  assign _T_1672 = $signed(_T_1671) & $signed(-33'sh10000000); 
  assign _T_1673 = $signed(_T_1672); 
  assign _T_1674 = $signed(_T_1673) == $signed(33'sh0); 
  assign _T_1676 = _T_1664 | _T_1669; 
  assign _T_1677 = _T_1676 | _T_1674; 
  assign _T_1808 = io_in_c_bits_opcode == 3'h4; 
  assign _T_1810 = _T_1677 | reset; 
  assign _T_1811 = _T_1810 == 1'h0; 
  assign _T_1813 = _T_1653 | reset; 
  assign _T_1814 = _T_1813 == 1'h0; 
  assign _T_1815 = io_in_c_bits_size >= 4'h3; 
  assign _T_1817 = _T_1815 | reset; 
  assign _T_1818 = _T_1817 == 1'h0; 
  assign _T_1820 = _T_1659 | reset; 
  assign _T_1821 = _T_1820 == 1'h0; 
  assign _T_1822 = io_in_c_bits_param <= 3'h5; 
  assign _T_1824 = _T_1822 | reset; 
  assign _T_1825 = _T_1824 == 1'h0; 
  assign _T_1826 = io_in_c_bits_corrupt == 1'h0; 
  assign _T_1828 = _T_1826 | reset; 
  assign _T_1829 = _T_1828 == 1'h0; 
  assign _T_1830 = io_in_c_bits_opcode == 3'h5; 
  assign _T_1848 = io_in_c_bits_opcode == 3'h6; 
  assign _T_1863 = io_in_c_bits_size <= 4'h6; 
  assign _T_1871 = _T_1863 & _T_1674; 
  assign _T_1875 = _T_1871 | reset; 
  assign _T_1876 = _T_1875 == 1'h0; 
  assign _T_1945 = _T_1585 ? _T_1863 : 1'h0; 
  assign _T_1962 = _T_1945 | reset; 
  assign _T_1963 = _T_1962 == 1'h0; 
  assign _T_1974 = io_in_c_bits_param <= 3'h2; 
  assign _T_1976 = _T_1974 | reset; 
  assign _T_1977 = _T_1976 == 1'h0; 
  assign _T_1982 = io_in_c_bits_opcode == 3'h7; 
  assign _T_2112 = io_in_c_bits_opcode == 3'h0; 
  assign _T_2122 = io_in_c_bits_param == 3'h0; 
  assign _T_2124 = _T_2122 | reset; 
  assign _T_2125 = _T_2124 == 1'h0; 
  assign _T_2130 = io_in_c_bits_opcode == 3'h1; 
  assign _T_2144 = io_in_c_bits_opcode == 3'h2; 
  assign _T_2162 = io_in_e_bits_sink < 1'h1; 
  assign _T_2164 = _T_2162 | reset; 
  assign _T_2165 = _T_2164 == 1'h0; 
  assign _T_2166 = io_in_a_ready & io_in_a_valid; 
  assign _T_2171 = _T_80[7:3]; 
  assign _T_2172 = io_in_a_bits_opcode[2]; 
  assign _T_2173 = _T_2172 == 1'h0; 
  assign _T_2177 = _T_2175 - 5'h1; 
  assign _T_2178 = _T_2175 == 5'h0; 
  assign _T_2191 = _T_2178 == 1'h0; 
  assign _T_2192 = io_in_a_valid & _T_2191; 
  assign _T_2193 = io_in_a_bits_opcode == _T_2186; 
  assign _T_2195 = _T_2193 | reset; 
  assign _T_2196 = _T_2195 == 1'h0; 
  assign _T_2197 = io_in_a_bits_param == _T_2187; 
  assign _T_2199 = _T_2197 | reset; 
  assign _T_2200 = _T_2199 == 1'h0; 
  assign _T_2201 = io_in_a_bits_size == _T_2188; 
  assign _T_2203 = _T_2201 | reset; 
  assign _T_2204 = _T_2203 == 1'h0; 
  assign _T_2205 = io_in_a_bits_source == _T_2189; 
  assign _T_2207 = _T_2205 | reset; 
  assign _T_2208 = _T_2207 == 1'h0; 
  assign _T_2209 = io_in_a_bits_address == _T_2190; 
  assign _T_2211 = _T_2209 | reset; 
  assign _T_2212 = _T_2211 == 1'h0; 
  assign _T_2214 = _T_2166 & _T_2178; 
  assign _T_2215 = io_in_d_ready & io_in_d_valid; 
  assign _T_2217 = 23'hff << io_in_d_bits_size; 
  assign _T_2218 = _T_2217[7:0]; 
  assign _T_2219 = ~ _T_2218; 
  assign _T_2220 = _T_2219[7:3]; 
  assign _T_2221 = io_in_d_bits_opcode[0]; 
  assign _T_2225 = _T_2223 - 5'h1; 
  assign _T_2226 = _T_2223 == 5'h0; 
  assign _T_2240 = _T_2226 == 1'h0; 
  assign _T_2241 = io_in_d_valid & _T_2240; 
  assign _T_2242 = io_in_d_bits_opcode == _T_2234; 
  assign _T_2244 = _T_2242 | reset; 
  assign _T_2245 = _T_2244 == 1'h0; 
  assign _T_2246 = io_in_d_bits_param == _T_2235; 
  assign _T_2248 = _T_2246 | reset; 
  assign _T_2249 = _T_2248 == 1'h0; 
  assign _T_2250 = io_in_d_bits_size == _T_2236; 
  assign _T_2252 = _T_2250 | reset; 
  assign _T_2253 = _T_2252 == 1'h0; 
  assign _T_2254 = io_in_d_bits_source == _T_2237; 
  assign _T_2256 = _T_2254 | reset; 
  assign _T_2257 = _T_2256 == 1'h0; 
  assign _T_2258 = io_in_d_bits_sink == _T_2238; 
  assign _T_2260 = _T_2258 | reset; 
  assign _T_2261 = _T_2260 == 1'h0; 
  assign _T_2262 = io_in_d_bits_denied == _T_2239; 
  assign _T_2264 = _T_2262 | reset; 
  assign _T_2265 = _T_2264 == 1'h0; 
  assign _T_2267 = _T_2215 & _T_2226; 
  assign _T_2317 = io_in_c_ready & io_in_c_valid; 
  assign _T_2322 = _T_1657[7:3]; 
  assign _T_2323 = io_in_c_bits_opcode[0]; 
  assign _T_2327 = _T_2325 - 5'h1; 
  assign _T_2328 = _T_2325 == 5'h0; 
  assign _T_2341 = _T_2328 == 1'h0; 
  assign _T_2342 = io_in_c_valid & _T_2341; 
  assign _T_2343 = io_in_c_bits_opcode == _T_2336; 
  assign _T_2345 = _T_2343 | reset; 
  assign _T_2346 = _T_2345 == 1'h0; 
  assign _T_2347 = io_in_c_bits_param == _T_2337; 
  assign _T_2349 = _T_2347 | reset; 
  assign _T_2350 = _T_2349 == 1'h0; 
  assign _T_2351 = io_in_c_bits_size == _T_2338; 
  assign _T_2353 = _T_2351 | reset; 
  assign _T_2354 = _T_2353 == 1'h0; 
  assign _T_2355 = io_in_c_bits_source == _T_2339; 
  assign _T_2357 = _T_2355 | reset; 
  assign _T_2358 = _T_2357 == 1'h0; 
  assign _T_2359 = io_in_c_bits_address == _T_2340; 
  assign _T_2361 = _T_2359 | reset; 
  assign _T_2362 = _T_2361 == 1'h0; 
  assign _T_2364 = _T_2317 & _T_2328; 
  assign _T_2377 = _T_2375 - 5'h1; 
  assign _T_2378 = _T_2375 == 5'h0; 
  assign _T_2396 = _T_2394 - 5'h1; 
  assign _T_2397 = _T_2394 == 5'h0; 
  assign _T_2407 = _T_2166 & _T_2378; 
  assign _T_2409 = 128'h1 << io_in_a_bits_source; 
  assign _T_2410 = _T_2365 >> io_in_a_bits_source; 
  assign _T_2411 = _T_2410[0]; 
  assign _T_2412 = _T_2411 == 1'h0; 
  assign _T_2414 = _T_2412 | reset; 
  assign _T_2415 = _T_2414 == 1'h0; 
  assign _GEN_27 = _T_2407 ? _T_2409 : 128'h0; 
  assign _T_2419 = _T_2215 & _T_2397; 
  assign _T_2421 = _T_904 == 1'h0; 
  assign _T_2422 = _T_2419 & _T_2421; 
  assign _T_2423 = 128'h1 << io_in_d_bits_source; 
  assign _T_2424 = _GEN_27 | _T_2365; 
  assign _T_2425 = _T_2424 >> io_in_d_bits_source; 
  assign _T_2426 = _T_2425[0]; 
  assign _T_2428 = _T_2426 | reset; 
  assign _T_2429 = _T_2428 == 1'h0; 
  assign _GEN_28 = _T_2422 ? _T_2423 : 128'h0; 
  assign _T_2430 = _GEN_27 != _GEN_28; 
  assign _T_2431 = _GEN_27 != 128'h0; 
  assign _T_2432 = _T_2431 == 1'h0; 
  assign _T_2433 = _T_2430 | _T_2432; 
  assign _T_2435 = _T_2433 | reset; 
  assign _T_2436 = _T_2435 == 1'h0; 
  assign _T_2437 = _T_2365 | _GEN_27; 
  assign _T_2438 = ~ _GEN_28; 
  assign _T_2439 = _T_2437 & _T_2438; 
  assign _T_2441 = _T_2365 != 128'h0; 
  assign _T_2442 = _T_2441 == 1'h0; 
  assign _T_2443 = plusarg_reader_out == 32'h0; 
  assign _T_2444 = _T_2442 | _T_2443; 
  assign _T_2445 = _T_2440 < plusarg_reader_out; 
  assign _T_2446 = _T_2444 | _T_2445; 
  assign _T_2448 = _T_2446 | reset; 
  assign _T_2449 = _T_2448 == 1'h0; 
  assign _T_2451 = _T_2440 + 32'h1; 
  assign _T_2454 = _T_2166 | _T_2215; 
  assign _T_2466 = _T_2464 - 5'h1; 
  assign _T_2467 = _T_2464 == 5'h0; 
  assign _T_2477 = _T_2215 & _T_2467; 
  assign _T_2478 = io_in_d_bits_opcode[2]; 
  assign _T_2479 = io_in_d_bits_opcode[1]; 
  assign _T_2480 = _T_2479 == 1'h0; 
  assign _T_2481 = _T_2478 & _T_2480; 
  assign _T_2482 = _T_2477 & _T_2481; 
  assign _T_2483 = 2'h1 << io_in_d_bits_sink; 
  assign _T_2484 = _T_2455 >> io_in_d_bits_sink; 
  assign _T_2486 = _T_2484 == 1'h0; 
  assign _T_2488 = _T_2486 | reset; 
  assign _T_2489 = _T_2488 == 1'h0; 
  assign _GEN_31 = _T_2482 ? _T_2483 : 2'h0; 
  assign _T_2491 = io_in_e_ready & io_in_e_valid; 
  assign _T_2494 = 2'h1 << io_in_e_bits_sink; 
  assign _T_2475 = _GEN_31[0]; 
  assign _T_2495 = _T_2475 | _T_2455; 
  assign _T_2496 = _T_2495 >> io_in_e_bits_sink; 
  assign _T_2499 = _T_2496 | reset; 
  assign _T_2500 = _T_2499 == 1'h0; 
  assign _GEN_32 = _T_2491 ? _T_2494 : 2'h0; 
  assign _T_2501 = _T_2455 | _T_2475; 
  assign _T_2490 = _GEN_32[0]; 
  assign _T_2502 = ~ _T_2490; 
  assign _T_2503 = _T_2501 & _T_2502; 
  assign _GEN_35 = io_in_a_valid & _T_277; 
  assign _GEN_51 = io_in_a_valid & _T_416; 
  assign _GEN_69 = io_in_a_valid & _T_559; 
  assign _GEN_81 = io_in_a_valid & _T_604; 
  assign _GEN_91 = io_in_a_valid & _T_650; 
  assign _GEN_101 = io_in_a_valid & _T_698; 
  assign _GEN_111 = io_in_a_valid & _T_741; 
  assign _GEN_121 = io_in_a_valid & _T_784; 
  assign _GEN_131 = io_in_d_valid & _T_904; 
  assign _GEN_141 = io_in_d_valid & _T_924; 
  assign _GEN_153 = io_in_d_valid & _T_952; 
  assign _GEN_165 = io_in_d_valid & _T_981; 
  assign _GEN_171 = io_in_d_valid & _T_998; 
  assign _GEN_177 = io_in_d_valid & _T_1016; 
  assign _GEN_183 = io_in_c_valid & _T_1808; 
  assign _GEN_195 = io_in_c_valid & _T_1830; 
  assign _GEN_205 = io_in_c_valid & _T_1848; 
  assign _GEN_219 = io_in_c_valid & _T_1982; 
  assign _GEN_231 = io_in_c_valid & _T_2112; 
  assign _GEN_241 = io_in_c_valid & _T_2130; 
  assign _GEN_249 = io_in_c_valid & _T_2144; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2175 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_2186 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2187 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_2188 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_2189 = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_2190 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_2223 = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_2234 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_2235 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_2236 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_2237 = _RAND_10[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_2238 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_2239 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_2325 = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_2336 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_2337 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_2338 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_2339 = _RAND_17[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_2340 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {4{`RANDOM}};
  _T_2365 = _RAND_19[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_2375 = _RAND_20[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_2394 = _RAND_21[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_2440 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_2455 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_2464 = _RAND_24[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_2175 <= 5'h0;
    end else begin
      if (_T_2166) begin
        if (_T_2178) begin
          if (_T_2173) begin
            _T_2175 <= _T_2171;
          end else begin
            _T_2175 <= 5'h0;
          end
        end else begin
          _T_2175 <= _T_2177;
        end
      end
    end
    if (_T_2214) begin
      _T_2186 <= io_in_a_bits_opcode;
    end
    if (_T_2214) begin
      _T_2187 <= io_in_a_bits_param;
    end
    if (_T_2214) begin
      _T_2188 <= io_in_a_bits_size;
    end
    if (_T_2214) begin
      _T_2189 <= io_in_a_bits_source;
    end
    if (_T_2214) begin
      _T_2190 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_2223 <= 5'h0;
    end else begin
      if (_T_2215) begin
        if (_T_2226) begin
          if (_T_2221) begin
            _T_2223 <= _T_2220;
          end else begin
            _T_2223 <= 5'h0;
          end
        end else begin
          _T_2223 <= _T_2225;
        end
      end
    end
    if (_T_2267) begin
      _T_2234 <= io_in_d_bits_opcode;
    end
    if (_T_2267) begin
      _T_2235 <= io_in_d_bits_param;
    end
    if (_T_2267) begin
      _T_2236 <= io_in_d_bits_size;
    end
    if (_T_2267) begin
      _T_2237 <= io_in_d_bits_source;
    end
    if (_T_2267) begin
      _T_2238 <= io_in_d_bits_sink;
    end
    if (_T_2267) begin
      _T_2239 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_2325 <= 5'h0;
    end else begin
      if (_T_2317) begin
        if (_T_2328) begin
          if (_T_2323) begin
            _T_2325 <= _T_2322;
          end else begin
            _T_2325 <= 5'h0;
          end
        end else begin
          _T_2325 <= _T_2327;
        end
      end
    end
    if (_T_2364) begin
      _T_2336 <= io_in_c_bits_opcode;
    end
    if (_T_2364) begin
      _T_2337 <= io_in_c_bits_param;
    end
    if (_T_2364) begin
      _T_2338 <= io_in_c_bits_size;
    end
    if (_T_2364) begin
      _T_2339 <= io_in_c_bits_source;
    end
    if (_T_2364) begin
      _T_2340 <= io_in_c_bits_address;
    end
    if (reset) begin
      _T_2365 <= 128'h0;
    end else begin
      _T_2365 <= _T_2439;
    end
    if (reset) begin
      _T_2375 <= 5'h0;
    end else begin
      if (_T_2166) begin
        if (_T_2378) begin
          if (_T_2173) begin
            _T_2375 <= _T_2171;
          end else begin
            _T_2375 <= 5'h0;
          end
        end else begin
          _T_2375 <= _T_2377;
        end
      end
    end
    if (reset) begin
      _T_2394 <= 5'h0;
    end else begin
      if (_T_2215) begin
        if (_T_2397) begin
          if (_T_2221) begin
            _T_2394 <= _T_2220;
          end else begin
            _T_2394 <= 5'h0;
          end
        end else begin
          _T_2394 <= _T_2396;
        end
      end
    end
    if (reset) begin
      _T_2440 <= 32'h0;
    end else begin
      if (_T_2454) begin
        _T_2440 <= 32'h0;
      end else begin
        _T_2440 <= _T_2451;
      end
    end
    if (reset) begin
      _T_2455 <= 1'h0;
    end else begin
      _T_2455 <= _T_2503;
    end
    if (reset) begin
      _T_2464 <= 5'h0;
    end else begin
      if (_T_2215) begin
        if (_T_2467) begin
          if (_T_2221) begin
            _T_2464 <= _T_2220;
          end else begin
            _T_2464 <= 5'h0;
          end
        end else begin
          _T_2464 <= _T_2466;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel has invalid opcode (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:39 assert (TLMessages.isA(bundle.opcode), \"'A' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:46 assert (visible(edge.address(bundle), bundle.source, edge), \"'A' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_305) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:49 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_305) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_392) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:50 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_392) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:51 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_399) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:52 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_399) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:53 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_406) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:54 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_406) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_411) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:55 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_411) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_35 & _T_415) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:56 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_35 & _T_415) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_305) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:60 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_305) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_392) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:61 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_392) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:62 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_399) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:63 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_399) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:64 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_406) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:65 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_406) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_549) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:66 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_549) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_411) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:67 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_411) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_51 & _T_415) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:68 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_51 & _T_415) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_585) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:72 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & _T_585) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:73 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:74 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_595) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:75 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & _T_595) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:76 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & _T_599) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_415) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:77 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_69 & _T_415) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_81 & _T_635) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:81 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_81 & _T_635) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_81 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_81 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_81 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_81 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_81 & _T_595) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_81 & _T_595) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_81 & _T_599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:85 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_81 & _T_599) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_635) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:89 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_635) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_595) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:92 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_595) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_697) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:93 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_697) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_305) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:97 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_305) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_736) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:100 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_736) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_599) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & _T_305) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:105 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & _T_305) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & _T_779) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:108 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & _T_779) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & _T_599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:109 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & _T_599) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_305) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:113 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_305) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_395) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:114 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_395) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_402) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:115 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_402) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_599) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:116 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_599) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_415) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:117 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_415) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_830) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:268 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_830) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_907) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:276 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_907) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_911) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:277 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_911) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_915) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:278 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_915) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_919) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:279 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_919) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_131 & _T_923) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:280 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_131 & _T_923) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_907) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:284 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_907) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_930) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:285 assert (sink_ok, \"'D' channel Grant carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_930) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_911) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:286 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_911) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_938) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:287 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_938) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_942) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:288 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_942) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_919) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:289 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_919) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is denied (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:290 assert (deny_put_ok || !bundle.denied, \"'D' channel Grant is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_907) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:294 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_907) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_930) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:295 assert (sink_ok, \"'D' channel GrantData carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_930) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_911) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:296 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_911) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_938) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:297 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_938) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_942) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:298 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_942) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_975) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:299 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_975) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:300 assert (deny_get_ok || !bundle.denied, \"'D' channel GrantData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & _T_907) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:304 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & _T_907) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & _T_915) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:306 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & _T_915) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_165 & _T_919) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:307 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_165 & _T_919) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is denied (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:308 assert (deny_put_ok || !bundle.denied, \"'D' channel AccessAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_907) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:312 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_907) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_915) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:314 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_915) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_975) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:315 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_975) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:316 assert (deny_get_ok || !bundle.denied, \"'D' channel AccessAckData is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_177 & _T_907) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:320 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_177 & _T_907) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_177 & _T_915) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:322 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_177 & _T_915) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_177 & _T_919) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:323 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_177 & _T_919) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is denied (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:324 assert (deny_put_ok || !bundle.denied, \"'D' channel HintAck is denied\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel has invalid opcode (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:122 assert (TLMessages.isB(bundle.opcode), \"'B' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:124 assert (visible(edge.address(bundle), bundle.source, edge), \"'B' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Probe type unsupported by client (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:133 assert (edge.client.supportsProbe(bundle.source, bundle.size), \"'B' channel carries Probe type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:134 assert (address_ok, \"'B' channel Probe carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries source that is not first source (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:135 assert (legal_source, \"'B' channel Probe carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:136 assert (is_aligned, \"'B' channel Probe address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:137 assert (TLPermissions.isCap(bundle.param), \"'B' channel Probe carries invalid cap param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe contains invalid mask (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:138 assert (bundle.mask === mask, \"'B' channel Probe contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe is corrupt (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:139 assert (!bundle.corrupt, \"'B' channel Probe is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Get type unsupported by client (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:143 assert (edge.client.supportsGet(bundle.source, bundle.size), \"'B' channel carries Get type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries unmanaged address (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:144 assert (address_ok, \"'B' channel Get carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries source that is not first source (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:145 assert (legal_source, \"'B' channel Get carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:146 assert (is_aligned, \"'B' channel Get address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries invalid param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:147 assert (bundle.param === UInt(0), \"'B' channel Get carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get contains invalid mask (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:148 assert (bundle.mask === mask, \"'B' channel Get contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get is corrupt (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:149 assert (!bundle.corrupt, \"'B' channel Get is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutFull type unsupported by client (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:153 assert (edge.client.supportsPutFull(bundle.source, bundle.size), \"'B' channel carries PutFull type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries unmanaged address (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:154 assert (address_ok, \"'B' channel PutFull carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries source that is not first source (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:155 assert (legal_source, \"'B' channel PutFull carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:156 assert (is_aligned, \"'B' channel PutFull address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries invalid param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:157 assert (bundle.param === UInt(0), \"'B' channel PutFull carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull contains invalid mask (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:158 assert (bundle.mask === mask, \"'B' channel PutFull contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutPartial type unsupported by client (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:162 assert (edge.client.supportsPutPartial(bundle.source, bundle.size), \"'B' channel carries PutPartial type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:163 assert (address_ok, \"'B' channel PutPartial carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:164 assert (legal_source, \"'B' channel PutPartial carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:165 assert (is_aligned, \"'B' channel PutPartial address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries invalid param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:166 assert (bundle.param === UInt(0), \"'B' channel PutPartial carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial contains invalid mask (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:167 assert ((bundle.mask & ~mask) === UInt(0), \"'B' channel PutPartial contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Arithmetic type unsupported by client (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:171 assert (edge.client.supportsArithmetic(bundle.source, bundle.size), \"'B' channel carries Arithmetic type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:172 assert (address_ok, \"'B' channel Arithmetic carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:173 assert (legal_source, \"'B' channel Arithmetic carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:174 assert (is_aligned, \"'B' channel Arithmetic address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries invalid opcode param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:175 assert (TLAtomics.isArithmetic(bundle.param), \"'B' channel Arithmetic carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:176 assert (bundle.mask === mask, \"'B' channel Arithmetic contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Logical type unsupported by client (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:180 assert (edge.client.supportsLogical(bundle.source, bundle.size), \"'B' channel carries Logical type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries unmanaged address (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:181 assert (address_ok, \"'B' channel Logical carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries source that is not first source (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:182 assert (legal_source, \"'B' channel Logical carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:183 assert (is_aligned, \"'B' channel Logical address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries invalid opcode param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:184 assert (TLAtomics.isLogical(bundle.param), \"'B' channel Logical carries invalid opcode param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical contains invalid mask (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:185 assert (bundle.mask === mask, \"'B' channel Logical contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Hint type unsupported by client (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:189 assert (edge.client.supportsHint(bundle.source, bundle.size), \"'B' channel carries Hint type unsupported by client\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries unmanaged address (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:190 assert (address_ok, \"'B' channel Hint carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries source that is not first source (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:191 assert (legal_source, \"'B' channel Hint carries source that is not first source\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:192 assert (is_aligned, \"'B' channel Hint address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint contains invalid mask (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:193 assert (bundle.mask === mask, \"'B' channel Hint contains invalid mask\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint is corrupt (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:194 assert (!bundle.corrupt, \"'B' channel Hint is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel has invalid opcode (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:199 assert (TLMessages.isC(bundle.opcode), \"'C' channel has invalid opcode\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:205 assert (visible(edge.address(bundle), bundle.source, edge), \"'C' channel carries an address illegal for the specified bank visibility\")\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_1811) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:208 assert (address_ok, \"'C' channel ProbeAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_1811) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_1814) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:209 assert (source_ok, \"'C' channel ProbeAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_1814) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_1818) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:210 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAck smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_1818) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_1821) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:211 assert (is_aligned, \"'C' channel ProbeAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_1821) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_1825) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:212 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAck carries invalid report param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_1825) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & _T_1829) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck is corrupt (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:213 assert (!bundle.corrupt, \"'C' channel ProbeAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & _T_1829) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1811) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:217 assert (address_ok, \"'C' channel ProbeAckData carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1811) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1814) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:218 assert (source_ok, \"'C' channel ProbeAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1814) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1818) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:219 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ProbeAckData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1818) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1821) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:220 assert (is_aligned, \"'C' channel ProbeAckData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1821) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_1825) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:221 assert (TLPermissions.isReport(bundle.param), \"'C' channel ProbeAckData carries invalid report param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_1825) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1876) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:225 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries Release type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1876) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1963) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:226 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1963) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1814) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:227 assert (source_ok, \"'C' channel Release carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1814) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1818) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:228 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel Release smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1818) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1821) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:229 assert (is_aligned, \"'C' channel Release address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1821) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1977) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid shrink param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:230 assert (TLPermissions.isShrink(bundle.param), \"'C' channel Release carries invalid shrink param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1977) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_1829) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release is corrupt (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:231 assert (!bundle.corrupt, \"'C' channel Release is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_1829) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1876) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:235 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'C' channel carries ReleaseData type unsupported by manager\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1876) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1963) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:236 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'C' channel carries Release from a client which does not support Probe\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1963) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1814) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:237 assert (source_ok, \"'C' channel ReleaseData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1814) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1818) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:238 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'C' channel ReleaseData smaller than a beat\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1818) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1821) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:239 assert (is_aligned, \"'C' channel ReleaseData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1821) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_219 & _T_1977) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid shrink param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:240 assert (TLPermissions.isShrink(bundle.param), \"'C' channel ReleaseData carries invalid shrink param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_219 & _T_1977) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1811) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:244 assert (address_ok, \"'C' channel AccessAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1811) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1814) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:245 assert (source_ok, \"'C' channel AccessAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1814) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1821) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:246 assert (is_aligned, \"'C' channel AccessAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1821) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_2125) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:247 assert (bundle.param === UInt(0), \"'C' channel AccessAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_2125) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_231 & _T_1829) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck is corrupt (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:248 assert (!bundle.corrupt, \"'C' channel AccessAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_231 & _T_1829) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1811) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:252 assert (address_ok, \"'C' channel AccessAckData carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1811) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1814) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:253 assert (source_ok, \"'C' channel AccessAckData carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1814) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1821) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:254 assert (is_aligned, \"'C' channel AccessAckData address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1821) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_2125) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:255 assert (bundle.param === UInt(0), \"'C' channel AccessAckData carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_2125) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_249 & _T_1811) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:259 assert (address_ok, \"'C' channel HintAck carries unmanaged address\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_249 & _T_1811) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_249 & _T_1814) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:260 assert (source_ok, \"'C' channel HintAck carries invalid source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_249 & _T_1814) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_249 & _T_1821) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:261 assert (is_aligned, \"'C' channel HintAck address not aligned to size\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_249 & _T_1821) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_249 & _T_2125) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:262 assert (bundle.param === UInt(0), \"'C' channel HintAck carries invalid param\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_249 & _T_2125) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_249 & _T_1829) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck is corrupt (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:263 assert (!bundle.corrupt, \"'C' channel HintAck is corrupt\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_249 & _T_1829) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_e_valid & _T_2165) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channels carries invalid sink ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:330 assert (sink_ok, \"'E' channels carries invalid sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_e_valid & _T_2165) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2192 & _T_2196) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:355 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2192 & _T_2196) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2192 & _T_2200) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:356 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2192 & _T_2200) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2192 & _T_2204) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:357 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2192 & _T_2204) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2192 & _T_2208) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:358 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2192 & _T_2208) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2192 & _T_2212) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:359 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2192 & _T_2212) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2241 & _T_2245) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:425 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2241 & _T_2245) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2241 & _T_2249) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:426 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2241 & _T_2249) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2241 & _T_2253) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:427 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2241 & _T_2253) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2241 & _T_2257) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:428 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2241 & _T_2257) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2241 & _T_2261) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:429 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2241 & _T_2261) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2241 & _T_2265) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:430 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2241 & _T_2265) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:378 assert (b.bits.opcode === opcode, \"'B' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:379 assert (b.bits.param  === param,  \"'B' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel size changed within multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:380 assert (b.bits.size   === size,   \"'B' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel source changed within multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:381 assert (b.bits.source === source, \"'B' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:382 assert (b.bits.address=== address,\"'B' channel addresss changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2342 & _T_2346) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:401 assert (c.bits.opcode === opcode, \"'C' channel opcode changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2342 & _T_2346) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2342 & _T_2350) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:402 assert (c.bits.param  === param,  \"'C' channel param changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2342 & _T_2350) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2342 & _T_2354) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:403 assert (c.bits.size   === size,   \"'C' channel size changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2342 & _T_2354) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2342 & _T_2358) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:404 assert (c.bits.source === source, \"'C' channel source changed within multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2342 & _T_2358) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2342 & _T_2362) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:405 assert (c.bits.address=== address,\"'C' channel address changed with multibeat operation\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2342 & _T_2362) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2407 & _T_2415) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:460 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2407 & _T_2415) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2422 & _T_2429) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:467 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2422 & _T_2429) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2436) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:471 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2436) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2449) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:479 assert (!inflight.orR || limit === UInt(0) || watchdog < limit, \"TileLink timeout expired\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2449) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2482 & _T_2489) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:494 assert(!inflight(bundle.d.bits.sink), \"'D' channel re-used a sink ID\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2482 & _T_2489) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2491 & _T_2500) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at ChiplinkTest.scala:362:8)\n    at Monitor.scala:500 assert((d_set | inflight)(bundle.e.bits.sink), \"'E' channel acknowledged for nothing inflight\" + extra)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2491 & _T_2500) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLToAXI4_1( 
  input         clock, 
  input         reset, 
  output        auto_in_a_ready, 
  input         auto_in_a_valid, 
  input  [2:0]  auto_in_a_bits_opcode, 
  input  [2:0]  auto_in_a_bits_param, 
  input  [3:0]  auto_in_a_bits_size, 
  input  [6:0]  auto_in_a_bits_source, 
  input  [30:0] auto_in_a_bits_address, 
  input  [7:0]  auto_in_a_bits_mask, 
  input  [63:0] auto_in_a_bits_data, 
  input         auto_in_a_bits_corrupt, 
  input         auto_in_d_ready, 
  output        auto_in_d_valid, 
  output [2:0]  auto_in_d_bits_opcode, 
  output [3:0]  auto_in_d_bits_size, 
  output [6:0]  auto_in_d_bits_source, 
  output        auto_in_d_bits_denied, 
  output [63:0] auto_in_d_bits_data, 
  output        auto_in_d_bits_corrupt, 
  input         auto_out_awready, 
  output        auto_out_awvalid, 
  output [4:0]  auto_out_awid, 
  output [30:0] auto_out_awaddr, 
  output [7:0]  auto_out_awlen, 
  output [2:0]  auto_out_awsize, 
  output [1:0]  auto_out_awburst, 
  output        auto_out_awlock, 
  output [3:0]  auto_out_awcache, 
  output [2:0]  auto_out_awprot, 
  output [3:0]  auto_out_awqos, 
  output [10:0] auto_out_awuser, 
  output [63:0] auto_out_awinstret, 
  input         auto_out_wready, 
  output        auto_out_wvalid, 
  output [63:0] auto_out_wdata, 
  output [7:0]  auto_out_wstrb, 
  output        auto_out_wlast, 
  output        auto_out_bready, 
  input         auto_out_bvalid, 
  input  [4:0]  auto_out_bid, 
  input  [1:0]  auto_out_bresp, 
  input  [10:0] auto_out_buser, 
  input         auto_out_arready, 
  output        auto_out_arvalid, 
  output [4:0]  auto_out_arid, 
  output [30:0] auto_out_araddr, 
  output [7:0]  auto_out_arlen, 
  output [2:0]  auto_out_arsize, 
  output [1:0]  auto_out_arburst, 
  output        auto_out_arlock, 
  output [3:0]  auto_out_arcache, 
  output [2:0]  auto_out_arprot, 
  output [3:0]  auto_out_arqos, 
  output [10:0] auto_out_aruser, 
  output [63:0] auto_out_arinstret, 
  output        auto_out_rready, 
  input         auto_out_rvalid, 
  input  [4:0]  auto_out_rid, 
  input  [63:0] auto_out_rdata, 
  input  [1:0]  auto_out_rresp, 
  input  [10:0] auto_out_ruser, 
  input         auto_out_rlast 
);
  wire  TLMonitor_clock; 
  wire  TLMonitor_reset; 
  wire  TLMonitor_io_in_a_ready; 
  wire  TLMonitor_io_in_a_valid; 
  wire [2:0] TLMonitor_io_in_a_bits_opcode; 
  wire [2:0] TLMonitor_io_in_a_bits_param; 
  wire [3:0] TLMonitor_io_in_a_bits_size; 
  wire [6:0] TLMonitor_io_in_a_bits_source; 
  wire [30:0] TLMonitor_io_in_a_bits_address; 
  wire [7:0] TLMonitor_io_in_a_bits_mask; 
  wire  TLMonitor_io_in_a_bits_corrupt; 
  wire  TLMonitor_io_in_d_ready; 
  wire  TLMonitor_io_in_d_valid; 
  wire [2:0] TLMonitor_io_in_d_bits_opcode; 
  wire [3:0] TLMonitor_io_in_d_bits_size; 
  wire [6:0] TLMonitor_io_in_d_bits_source; 
  wire  TLMonitor_io_in_d_bits_denied; 
  wire  TLMonitor_io_in_d_bits_corrupt; 
  wire  Queue_clock; 
  wire  Queue_reset; 
  wire  Queue_io_enq_ready; 
  wire  Queue_io_enq_valid; 
  wire [63:0] Queue_io_enq_bits_data; 
  wire [7:0] Queue_io_enq_bits_strb; 
  wire  Queue_io_enq_bits_last; 
  wire  Queue_io_deq_ready; 
  wire  Queue_io_deq_valid; 
  wire [63:0] Queue_io_deq_bits_data; 
  wire [7:0] Queue_io_deq_bits_strb; 
  wire  Queue_io_deq_bits_last; 
  wire  Queue_1_clock; 
  wire  Queue_1_reset; 
  wire  Queue_1_io_enq_ready; 
  wire  Queue_1_io_enq_valid; 
  wire [4:0] Queue_1_io_enq_bits_id; 
  wire [30:0] Queue_1_io_enq_bits_addr; 
  wire [7:0] Queue_1_io_enq_bits_len; 
  wire [2:0] Queue_1_io_enq_bits_size; 
  wire [10:0] Queue_1_io_enq_bits_user; 
  wire  Queue_1_io_enq_bits_wen; 
  wire  Queue_1_io_deq_ready; 
  wire  Queue_1_io_deq_valid; 
  wire [4:0] Queue_1_io_deq_bits_id; 
  wire [30:0] Queue_1_io_deq_bits_addr; 
  wire [7:0] Queue_1_io_deq_bits_len; 
  wire [2:0] Queue_1_io_deq_bits_size; 
  wire [1:0] Queue_1_io_deq_bits_burst; 
  wire  Queue_1_io_deq_bits_lock; 
  wire [3:0] Queue_1_io_deq_bits_cache; 
  wire [2:0] Queue_1_io_deq_bits_prot; 
  wire [3:0] Queue_1_io_deq_bits_qos; 
  wire [10:0] Queue_1_io_deq_bits_user; 
  wire [63:0] Queue_1_io_deq_bits_instret; 
  wire  Queue_1_io_deq_bits_wen; 
  wire  _T_12; 
  wire  _T_13; 
  reg [4:0] _T_330; 
  reg [31:0] _RAND_0;
  wire  _T_332; 
  wire  _T_355; 
  reg  _T_331; 
  reg [31:0] _RAND_1;
  wire  _T_354; 
  wire  _T_356; 
  wire  _T_357; 
  wire  _T_358; 
  reg [4:0] _T_301; 
  reg [31:0] _RAND_2;
  wire  _T_303; 
  wire  _T_326; 
  reg  _T_302; 
  reg [31:0] _RAND_3;
  wire  _T_325; 
  wire  _T_327; 
  wire  _T_328; 
  wire  _T_329; 
  reg [4:0] _T_272; 
  reg [31:0] _RAND_4;
  wire  _T_274; 
  wire  _T_297; 
  reg  _T_273; 
  reg [31:0] _RAND_5;
  wire  _T_296; 
  wire  _T_298; 
  wire  _T_299; 
  wire  _T_300; 
  reg [4:0] _T_243; 
  reg [31:0] _RAND_6;
  wire  _T_245; 
  wire  _T_268; 
  reg  _T_244; 
  reg [31:0] _RAND_7;
  wire  _T_267; 
  wire  _T_269; 
  wire  _T_270; 
  wire  _T_271; 
  reg [4:0] _T_214; 
  reg [31:0] _RAND_8;
  wire  _T_216; 
  wire  _T_239; 
  reg  _T_215; 
  reg [31:0] _RAND_9;
  wire  _T_238; 
  wire  _T_240; 
  wire  _T_241; 
  wire  _T_242; 
  reg [4:0] _T_185; 
  reg [31:0] _RAND_10;
  wire  _T_187; 
  wire  _T_210; 
  reg  _T_186; 
  reg [31:0] _RAND_11;
  wire  _T_209; 
  wire  _T_211; 
  wire  _T_212; 
  wire  _T_213; 
  reg [4:0] _T_156; 
  reg [31:0] _RAND_12;
  wire  _T_158; 
  wire  _T_181; 
  reg  _T_157; 
  reg [31:0] _RAND_13;
  wire  _T_180; 
  wire  _T_182; 
  wire  _T_183; 
  wire  _T_184; 
  reg  _T_779; 
  reg [31:0] _RAND_14;
  reg  _T_751; 
  reg [31:0] _RAND_15;
  reg  _T_723; 
  reg [31:0] _RAND_16;
  reg  _T_695; 
  reg [31:0] _RAND_17;
  reg  _T_667; 
  reg [31:0] _RAND_18;
  reg  _T_639; 
  reg [31:0] _RAND_19;
  reg  _T_611; 
  reg [31:0] _RAND_20;
  reg  _T_583; 
  reg [31:0] _RAND_21;
  reg  _T_555; 
  reg [31:0] _RAND_22;
  reg  _T_527; 
  reg [31:0] _RAND_23;
  reg  _T_499; 
  reg [31:0] _RAND_24;
  reg  _T_471; 
  reg [31:0] _RAND_25;
  reg  _T_443; 
  reg [31:0] _RAND_26;
  reg  _T_415; 
  reg [31:0] _RAND_27;
  reg  _T_387; 
  reg [31:0] _RAND_28;
  reg  _T_359; 
  reg [31:0] _RAND_29;
  wire  _GEN_131; 
  wire  _GEN_132; 
  wire  _GEN_133; 
  wire  _GEN_134; 
  wire  _GEN_135; 
  wire  _GEN_136; 
  wire  _GEN_137; 
  wire  _GEN_138; 
  wire  _GEN_139; 
  wire  _GEN_140; 
  wire  _GEN_141; 
  wire  _GEN_142; 
  wire  _GEN_143; 
  wire  _GEN_144; 
  wire  _GEN_145; 
  wire  _GEN_146; 
  wire  _GEN_147; 
  wire  _GEN_148; 
  wire  _GEN_149; 
  wire  _GEN_150; 
  wire  _GEN_151; 
  wire  _GEN_152; 
  wire  _GEN_153; 
  wire  _GEN_154; 
  wire  _GEN_155; 
  wire  _GEN_156; 
  wire  _GEN_157; 
  wire  _GEN_158; 
  wire  _GEN_159; 
  wire  _GEN_160; 
  wire  _GEN_161; 
  wire  _GEN_162; 
  wire  _GEN_163; 
  wire  _GEN_164; 
  wire  _GEN_165; 
  wire  _GEN_166; 
  wire  _GEN_167; 
  wire  _GEN_168; 
  wire  _GEN_169; 
  wire  _GEN_170; 
  wire  _GEN_171; 
  wire  _GEN_172; 
  wire  _GEN_173; 
  wire  _GEN_174; 
  wire  _GEN_175; 
  wire  _GEN_176; 
  wire  _GEN_177; 
  wire  _GEN_178; 
  wire  _GEN_179; 
  wire  _GEN_180; 
  wire  _GEN_181; 
  wire  _GEN_182; 
  wire  _GEN_183; 
  wire  _GEN_184; 
  wire  _GEN_185; 
  wire  _GEN_186; 
  wire  _GEN_187; 
  wire  _GEN_188; 
  wire  _GEN_189; 
  wire  _GEN_190; 
  wire  _GEN_191; 
  wire  _GEN_192; 
  wire  _GEN_193; 
  wire  _GEN_194; 
  wire  _GEN_195; 
  wire  _GEN_196; 
  wire  _GEN_197; 
  wire  _GEN_198; 
  wire  _GEN_199; 
  wire  _GEN_200; 
  wire  _GEN_201; 
  wire  _GEN_202; 
  wire  _GEN_203; 
  wire  _GEN_204; 
  wire  _GEN_205; 
  wire  _GEN_206; 
  wire  _GEN_207; 
  wire  _GEN_208; 
  wire  _GEN_209; 
  wire  _GEN_210; 
  wire  _GEN_211; 
  wire  _GEN_212; 
  wire  _GEN_213; 
  wire  _GEN_214; 
  wire  _GEN_215; 
  wire  _GEN_216; 
  wire  _GEN_217; 
  wire  _GEN_218; 
  wire  _GEN_219; 
  wire  _GEN_220; 
  wire  _GEN_221; 
  wire  _GEN_222; 
  wire  _GEN_223; 
  wire  _GEN_224; 
  wire  _GEN_225; 
  wire  _GEN_226; 
  wire  _GEN_227; 
  wire  _GEN_228; 
  wire  _GEN_229; 
  wire  _GEN_230; 
  wire  _GEN_231; 
  wire  _GEN_232; 
  wire  _GEN_233; 
  wire  _GEN_234; 
  wire  _GEN_235; 
  wire  _GEN_236; 
  wire  _GEN_237; 
  wire  _GEN_238; 
  wire  _GEN_239; 
  wire  _GEN_240; 
  wire  _GEN_241; 
  wire  _GEN_242; 
  wire  _GEN_243; 
  wire  _GEN_244; 
  wire  _GEN_245; 
  wire  _GEN_246; 
  wire  _GEN_247; 
  wire  _GEN_248; 
  wire  _GEN_249; 
  wire  _GEN_250; 
  wire  _GEN_251; 
  wire  _GEN_252; 
  wire  _GEN_253; 
  wire  _GEN_254; 
  wire  _GEN_255; 
  wire  _GEN_256; 
  wire  _GEN_257; 
  reg [4:0] _T_23; 
  reg [31:0] _RAND_30;
  wire  _T_26; 
  wire  _T_67; 
  wire  _T_68; 
  reg  _T_57; 
  reg [31:0] _RAND_31;
  wire  _T_49_ready; 
  wire  _T_69; 
  wire  _T_50_ready; 
  wire  _T_70; 
  wire  _T_71; 
  wire  _T_72; 
  wire  _T_14; 
  wire [22:0] _T_16; 
  wire [7:0] _T_17; 
  wire [7:0] _T_18; 
  wire [4:0] _T_19; 
  wire [4:0] _T_22; 
  wire [4:0] _T_25; 
  wire  _T_27; 
  wire  _T_28; 
  wire  _T_29; 
  wire [10:0] _T_43; 
  wire [10:0] _GEN_284; 
  wire [6:0] _T_45; 
  wire [3:0] _T_46; 
  wire [6:0] _T_47; 
  wire [3:0] _T_48; 
  wire  _T_52_bits_wen; 
  wire  _T_53; 
  wire  _T_52_valid; 
  wire  _T_59; 
  wire [4:0] _GEN_3; 
  wire [4:0] _GEN_4; 
  wire [4:0] _GEN_5; 
  wire [4:0] _GEN_6; 
  wire [4:0] _GEN_7; 
  wire [4:0] _GEN_8; 
  wire [4:0] _GEN_9; 
  wire [4:0] _GEN_10; 
  wire [4:0] _GEN_11; 
  wire [4:0] _GEN_12; 
  wire [4:0] _GEN_13; 
  wire [4:0] _GEN_14; 
  wire [4:0] _GEN_15; 
  wire [4:0] _GEN_16; 
  wire [4:0] _GEN_17; 
  wire [4:0] _GEN_18; 
  wire [4:0] _GEN_19; 
  wire [4:0] _GEN_20; 
  wire [4:0] _GEN_21; 
  wire [4:0] _GEN_22; 
  wire [4:0] _GEN_23; 
  wire [4:0] _GEN_24; 
  wire [4:0] _GEN_25; 
  wire [4:0] _GEN_26; 
  wire [4:0] _GEN_27; 
  wire [4:0] _GEN_28; 
  wire [4:0] _GEN_29; 
  wire [4:0] _GEN_30; 
  wire [4:0] _GEN_31; 
  wire [4:0] _GEN_32; 
  wire [4:0] _GEN_33; 
  wire [4:0] _GEN_34; 
  wire [4:0] _GEN_35; 
  wire [4:0] _GEN_36; 
  wire [4:0] _GEN_37; 
  wire [4:0] _GEN_38; 
  wire [4:0] _GEN_39; 
  wire [4:0] _GEN_40; 
  wire [4:0] _GEN_41; 
  wire [4:0] _GEN_42; 
  wire [4:0] _GEN_43; 
  wire [4:0] _GEN_44; 
  wire [4:0] _GEN_45; 
  wire [4:0] _GEN_46; 
  wire [4:0] _GEN_47; 
  wire [4:0] _GEN_48; 
  wire [4:0] _GEN_49; 
  wire [4:0] _GEN_50; 
  wire [4:0] _GEN_51; 
  wire [4:0] _GEN_52; 
  wire [4:0] _GEN_53; 
  wire [4:0] _GEN_54; 
  wire [4:0] _GEN_55; 
  wire [4:0] _GEN_56; 
  wire [4:0] _GEN_57; 
  wire [4:0] _GEN_58; 
  wire [4:0] _GEN_59; 
  wire [4:0] _GEN_60; 
  wire [4:0] _GEN_61; 
  wire [4:0] _GEN_62; 
  wire [4:0] _GEN_63; 
  wire [4:0] _GEN_64; 
  wire [4:0] _GEN_65; 
  wire [4:0] _GEN_66; 
  wire [4:0] _GEN_67; 
  wire [4:0] _GEN_68; 
  wire [4:0] _GEN_69; 
  wire [4:0] _GEN_70; 
  wire [4:0] _GEN_71; 
  wire [4:0] _GEN_72; 
  wire [4:0] _GEN_73; 
  wire [4:0] _GEN_74; 
  wire [4:0] _GEN_75; 
  wire [4:0] _GEN_76; 
  wire [4:0] _GEN_77; 
  wire [4:0] _GEN_78; 
  wire [4:0] _GEN_79; 
  wire [4:0] _GEN_80; 
  wire [4:0] _GEN_81; 
  wire [4:0] _GEN_82; 
  wire [4:0] _GEN_83; 
  wire [4:0] _GEN_84; 
  wire [4:0] _GEN_85; 
  wire [4:0] _GEN_86; 
  wire [4:0] _GEN_87; 
  wire [4:0] _GEN_88; 
  wire [4:0] _GEN_89; 
  wire [4:0] _GEN_90; 
  wire [4:0] _GEN_91; 
  wire [4:0] _GEN_92; 
  wire [4:0] _GEN_93; 
  wire [4:0] _GEN_94; 
  wire [4:0] _GEN_95; 
  wire [4:0] _GEN_96; 
  wire [4:0] _GEN_97; 
  wire [4:0] _GEN_98; 
  wire [4:0] _GEN_99; 
  wire [4:0] _GEN_100; 
  wire [4:0] _GEN_101; 
  wire [4:0] _GEN_102; 
  wire [4:0] _GEN_103; 
  wire [4:0] _GEN_104; 
  wire [4:0] _GEN_105; 
  wire [4:0] _GEN_106; 
  wire [4:0] _GEN_107; 
  wire [4:0] _GEN_108; 
  wire [4:0] _GEN_109; 
  wire [4:0] _GEN_110; 
  wire [4:0] _GEN_111; 
  wire [4:0] _GEN_112; 
  wire [4:0] _GEN_113; 
  wire [4:0] _GEN_114; 
  wire [4:0] _GEN_115; 
  wire [4:0] _GEN_116; 
  wire [4:0] _GEN_117; 
  wire [4:0] _GEN_118; 
  wire [4:0] _GEN_119; 
  wire [4:0] _GEN_120; 
  wire [4:0] _GEN_121; 
  wire [4:0] _GEN_122; 
  wire [4:0] _GEN_123; 
  wire [4:0] _GEN_124; 
  wire [4:0] _GEN_125; 
  wire [4:0] _GEN_126; 
  wire [4:0] _GEN_127; 
  wire [4:0] _GEN_128; 
  wire [4:0] _GEN_129; 
  wire [25:0] _T_61; 
  wire [10:0] _T_62; 
  wire [10:0] _T_63; 
  wire  _T_65; 
  wire [3:0] _T_66; 
  wire  _T_74; 
  wire  _T_75; 
  wire  _T_76; 
  wire  _T_77; 
  wire  _T_78; 
  wire  _T_81; 
  reg  _T_84; 
  reg [31:0] _RAND_32;
  wire  _T_85; 
  wire  _T_86; 
  wire  _T_87; 
  wire  _T_88; 
  wire  _T_90; 
  reg  _T_91; 
  reg [31:0] _RAND_33;
  wire  _T_93; 
  reg  _T_94; 
  reg [31:0] _RAND_34;
  wire  _GEN_260; 
  wire  _T_96; 
  wire  _T_97; 
  wire  _T_98; 
  wire [31:0] _T_103; 
  wire [22:0] _T_104; 
  wire  _T_105; 
  wire  _T_106; 
  wire  _T_107; 
  wire  _T_108; 
  wire  _T_109; 
  wire  _T_110; 
  wire  _T_111; 
  wire  _T_112; 
  wire  _T_113; 
  wire  _T_114; 
  wire  _T_115; 
  wire  _T_116; 
  wire  _T_117; 
  wire  _T_118; 
  wire  _T_119; 
  wire  _T_120; 
  wire  _T_121; 
  wire  _T_122; 
  wire  _T_123; 
  wire  _T_124; 
  wire  _T_125; 
  wire  _T_126; 
  wire  _T_127; 
  wire [4:0] _T_128; 
  wire [31:0] _T_130; 
  wire [22:0] _T_131; 
  wire  _T_132; 
  wire  _T_133; 
  wire  _T_134; 
  wire  _T_135; 
  wire  _T_136; 
  wire  _T_137; 
  wire  _T_138; 
  wire  _T_139; 
  wire  _T_140; 
  wire  _T_141; 
  wire  _T_142; 
  wire  _T_143; 
  wire  _T_144; 
  wire  _T_145; 
  wire  _T_146; 
  wire  _T_147; 
  wire  _T_148; 
  wire  _T_149; 
  wire  _T_150; 
  wire  _T_151; 
  wire  _T_152; 
  wire  _T_153; 
  wire  _T_154; 
  wire  _T_155; 
  wire  _T_159; 
  wire  _T_160; 
  wire  _T_161; 
  wire  _T_162; 
  wire  _T_163; 
  wire [4:0] _GEN_285; 
  wire [4:0] _T_165; 
  wire [4:0] _GEN_286; 
  wire [4:0] _T_167; 
  wire  _T_168; 
  wire  _T_169; 
  wire  _T_170; 
  wire  _T_172; 
  wire  _T_173; 
  wire  _T_174; 
  wire  _T_175; 
  wire  _T_176; 
  wire  _T_178; 
  wire  _T_179; 
  wire  _T_189; 
  wire  _T_190; 
  wire  _T_192; 
  wire [4:0] _GEN_287; 
  wire [4:0] _T_194; 
  wire [4:0] _GEN_288; 
  wire [4:0] _T_196; 
  wire  _T_197; 
  wire  _T_198; 
  wire  _T_199; 
  wire  _T_201; 
  wire  _T_202; 
  wire  _T_203; 
  wire  _T_204; 
  wire  _T_205; 
  wire  _T_207; 
  wire  _T_208; 
  wire  _T_218; 
  wire  _T_219; 
  wire  _T_221; 
  wire [4:0] _GEN_289; 
  wire [4:0] _T_223; 
  wire [4:0] _GEN_290; 
  wire [4:0] _T_225; 
  wire  _T_226; 
  wire  _T_227; 
  wire  _T_228; 
  wire  _T_230; 
  wire  _T_231; 
  wire  _T_232; 
  wire  _T_233; 
  wire  _T_234; 
  wire  _T_236; 
  wire  _T_237; 
  wire  _T_247; 
  wire  _T_248; 
  wire  _T_250; 
  wire [4:0] _GEN_291; 
  wire [4:0] _T_252; 
  wire [4:0] _GEN_292; 
  wire [4:0] _T_254; 
  wire  _T_255; 
  wire  _T_256; 
  wire  _T_257; 
  wire  _T_259; 
  wire  _T_260; 
  wire  _T_261; 
  wire  _T_262; 
  wire  _T_263; 
  wire  _T_265; 
  wire  _T_266; 
  wire  _T_276; 
  wire  _T_277; 
  wire  _T_279; 
  wire [4:0] _GEN_293; 
  wire [4:0] _T_281; 
  wire [4:0] _GEN_294; 
  wire [4:0] _T_283; 
  wire  _T_284; 
  wire  _T_285; 
  wire  _T_286; 
  wire  _T_288; 
  wire  _T_289; 
  wire  _T_290; 
  wire  _T_291; 
  wire  _T_292; 
  wire  _T_294; 
  wire  _T_295; 
  wire  _T_305; 
  wire  _T_306; 
  wire  _T_308; 
  wire [4:0] _GEN_295; 
  wire [4:0] _T_310; 
  wire [4:0] _GEN_296; 
  wire [4:0] _T_312; 
  wire  _T_313; 
  wire  _T_314; 
  wire  _T_315; 
  wire  _T_317; 
  wire  _T_318; 
  wire  _T_319; 
  wire  _T_320; 
  wire  _T_321; 
  wire  _T_323; 
  wire  _T_324; 
  wire  _T_334; 
  wire  _T_335; 
  wire  _T_337; 
  wire [4:0] _GEN_297; 
  wire [4:0] _T_339; 
  wire [4:0] _GEN_298; 
  wire [4:0] _T_341; 
  wire  _T_342; 
  wire  _T_343; 
  wire  _T_344; 
  wire  _T_346; 
  wire  _T_347; 
  wire  _T_348; 
  wire  _T_349; 
  wire  _T_350; 
  wire  _T_352; 
  wire  _T_353; 
  wire  _T_363; 
  wire  _T_364; 
  wire  _T_366; 
  wire  _T_368; 
  wire  _T_370; 
  wire  _T_371; 
  wire  _T_373; 
  wire  _T_375; 
  wire  _T_376; 
  wire  _T_377; 
  wire  _T_378; 
  wire  _T_379; 
  wire  _T_381; 
  wire  _T_382; 
  wire  _T_391; 
  wire  _T_392; 
  wire  _T_394; 
  wire  _T_396; 
  wire  _T_398; 
  wire  _T_399; 
  wire  _T_401; 
  wire  _T_403; 
  wire  _T_404; 
  wire  _T_405; 
  wire  _T_406; 
  wire  _T_407; 
  wire  _T_409; 
  wire  _T_410; 
  wire  _T_419; 
  wire  _T_420; 
  wire  _T_422; 
  wire  _T_424; 
  wire  _T_426; 
  wire  _T_427; 
  wire  _T_429; 
  wire  _T_431; 
  wire  _T_432; 
  wire  _T_433; 
  wire  _T_434; 
  wire  _T_435; 
  wire  _T_437; 
  wire  _T_438; 
  wire  _T_447; 
  wire  _T_448; 
  wire  _T_450; 
  wire  _T_452; 
  wire  _T_454; 
  wire  _T_455; 
  wire  _T_457; 
  wire  _T_459; 
  wire  _T_460; 
  wire  _T_461; 
  wire  _T_462; 
  wire  _T_463; 
  wire  _T_465; 
  wire  _T_466; 
  wire  _T_475; 
  wire  _T_476; 
  wire  _T_478; 
  wire  _T_480; 
  wire  _T_482; 
  wire  _T_483; 
  wire  _T_485; 
  wire  _T_487; 
  wire  _T_488; 
  wire  _T_489; 
  wire  _T_490; 
  wire  _T_491; 
  wire  _T_493; 
  wire  _T_494; 
  wire  _T_503; 
  wire  _T_504; 
  wire  _T_506; 
  wire  _T_508; 
  wire  _T_510; 
  wire  _T_511; 
  wire  _T_513; 
  wire  _T_515; 
  wire  _T_516; 
  wire  _T_517; 
  wire  _T_518; 
  wire  _T_519; 
  wire  _T_521; 
  wire  _T_522; 
  wire  _T_531; 
  wire  _T_532; 
  wire  _T_534; 
  wire  _T_536; 
  wire  _T_538; 
  wire  _T_539; 
  wire  _T_541; 
  wire  _T_543; 
  wire  _T_544; 
  wire  _T_545; 
  wire  _T_546; 
  wire  _T_547; 
  wire  _T_549; 
  wire  _T_550; 
  wire  _T_559; 
  wire  _T_560; 
  wire  _T_562; 
  wire  _T_564; 
  wire  _T_566; 
  wire  _T_567; 
  wire  _T_569; 
  wire  _T_571; 
  wire  _T_572; 
  wire  _T_573; 
  wire  _T_574; 
  wire  _T_575; 
  wire  _T_577; 
  wire  _T_578; 
  wire  _T_587; 
  wire  _T_588; 
  wire  _T_590; 
  wire  _T_592; 
  wire  _T_594; 
  wire  _T_595; 
  wire  _T_597; 
  wire  _T_599; 
  wire  _T_600; 
  wire  _T_601; 
  wire  _T_602; 
  wire  _T_603; 
  wire  _T_605; 
  wire  _T_606; 
  wire  _T_615; 
  wire  _T_616; 
  wire  _T_618; 
  wire  _T_620; 
  wire  _T_622; 
  wire  _T_623; 
  wire  _T_625; 
  wire  _T_627; 
  wire  _T_628; 
  wire  _T_629; 
  wire  _T_630; 
  wire  _T_631; 
  wire  _T_633; 
  wire  _T_634; 
  wire  _T_643; 
  wire  _T_644; 
  wire  _T_646; 
  wire  _T_648; 
  wire  _T_650; 
  wire  _T_651; 
  wire  _T_653; 
  wire  _T_655; 
  wire  _T_656; 
  wire  _T_657; 
  wire  _T_658; 
  wire  _T_659; 
  wire  _T_661; 
  wire  _T_662; 
  wire  _T_671; 
  wire  _T_672; 
  wire  _T_674; 
  wire  _T_676; 
  wire  _T_678; 
  wire  _T_679; 
  wire  _T_681; 
  wire  _T_683; 
  wire  _T_684; 
  wire  _T_685; 
  wire  _T_686; 
  wire  _T_687; 
  wire  _T_689; 
  wire  _T_690; 
  wire  _T_699; 
  wire  _T_700; 
  wire  _T_702; 
  wire  _T_704; 
  wire  _T_706; 
  wire  _T_707; 
  wire  _T_709; 
  wire  _T_711; 
  wire  _T_712; 
  wire  _T_713; 
  wire  _T_714; 
  wire  _T_715; 
  wire  _T_717; 
  wire  _T_718; 
  wire  _T_727; 
  wire  _T_728; 
  wire  _T_730; 
  wire  _T_732; 
  wire  _T_734; 
  wire  _T_735; 
  wire  _T_737; 
  wire  _T_739; 
  wire  _T_740; 
  wire  _T_741; 
  wire  _T_742; 
  wire  _T_743; 
  wire  _T_745; 
  wire  _T_746; 
  wire  _T_755; 
  wire  _T_756; 
  wire  _T_758; 
  wire  _T_760; 
  wire  _T_762; 
  wire  _T_763; 
  wire  _T_765; 
  wire  _T_767; 
  wire  _T_768; 
  wire  _T_769; 
  wire  _T_770; 
  wire  _T_771; 
  wire  _T_773; 
  wire  _T_774; 
  wire  _T_783; 
  wire  _T_784; 
  wire  _T_786; 
  wire  _T_788; 
  wire  _T_790; 
  wire  _T_791; 
  wire  _T_793; 
  wire  _T_795; 
  wire  _T_796; 
  wire  _T_797; 
  wire  _T_798; 
  wire  _T_799; 
  wire  _T_801; 
  wire  _T_802; 
  dual_TLMonitor_10 dual_TLMonitor ( 
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_io_in_a_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt)
  );
  dual_Queue_46 dual_Queue ( 
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_strb(Queue_io_enq_bits_strb),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_strb(Queue_io_deq_bits_strb),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  dual_Queue_57 Queue_1 ( 
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_id(Queue_1_io_enq_bits_id),
    .io_enq_bits_addr(Queue_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_user(Queue_1_io_enq_bits_user),
    .io_enq_bits_wen(Queue_1_io_enq_bits_wen),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_id(Queue_1_io_deq_bits_id),
    .io_deq_bits_addr(Queue_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_1_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_1_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_1_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_1_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_1_io_deq_bits_qos),
    .io_deq_bits_user(Queue_1_io_deq_bits_user),
    .io_deq_bits_instret(Queue_1_io_deq_bits_instret),
    .io_deq_bits_wen(Queue_1_io_deq_bits_wen)
  );
  assign _T_12 = auto_in_a_bits_opcode[2]; 
  assign _T_13 = _T_12 == 1'h0; 
  assign _T_332 = _T_330 == 5'h0; 
  assign _T_355 = _T_332 == 1'h0; 
  assign _T_354 = _T_331 != _T_13; 
  assign _T_356 = _T_355 & _T_354; 
  assign _T_357 = _T_330 == 5'h10; 
  assign _T_358 = _T_356 | _T_357; 
  assign _T_303 = _T_301 == 5'h0; 
  assign _T_326 = _T_303 == 1'h0; 
  assign _T_325 = _T_302 != _T_13; 
  assign _T_327 = _T_326 & _T_325; 
  assign _T_328 = _T_301 == 5'h10; 
  assign _T_329 = _T_327 | _T_328; 
  assign _T_274 = _T_272 == 5'h0; 
  assign _T_297 = _T_274 == 1'h0; 
  assign _T_296 = _T_273 != _T_13; 
  assign _T_298 = _T_297 & _T_296; 
  assign _T_299 = _T_272 == 5'h10; 
  assign _T_300 = _T_298 | _T_299; 
  assign _T_245 = _T_243 == 5'h0; 
  assign _T_268 = _T_245 == 1'h0; 
  assign _T_267 = _T_244 != _T_13; 
  assign _T_269 = _T_268 & _T_267; 
  assign _T_270 = _T_243 == 5'h10; 
  assign _T_271 = _T_269 | _T_270; 
  assign _T_216 = _T_214 == 5'h0; 
  assign _T_239 = _T_216 == 1'h0; 
  assign _T_238 = _T_215 != _T_13; 
  assign _T_240 = _T_239 & _T_238; 
  assign _T_241 = _T_214 == 5'h10; 
  assign _T_242 = _T_240 | _T_241; 
  assign _T_187 = _T_185 == 5'h0; 
  assign _T_210 = _T_187 == 1'h0; 
  assign _T_209 = _T_186 != _T_13; 
  assign _T_211 = _T_210 & _T_209; 
  assign _T_212 = _T_185 == 5'h10; 
  assign _T_213 = _T_211 | _T_212; 
  assign _T_158 = _T_156 == 5'h0; 
  assign _T_181 = _T_158 == 1'h0; 
  assign _T_180 = _T_157 != _T_13; 
  assign _T_182 = _T_181 & _T_180; 
  assign _T_183 = _T_156 == 5'h10; 
  assign _T_184 = _T_182 | _T_183; 
  assign _GEN_131 = 7'h1 == auto_in_a_bits_source ? _T_387 : _T_359; 
  assign _GEN_132 = 7'h2 == auto_in_a_bits_source ? _T_415 : _GEN_131; 
  assign _GEN_133 = 7'h3 == auto_in_a_bits_source ? _T_443 : _GEN_132; 
  assign _GEN_134 = 7'h4 == auto_in_a_bits_source ? _T_471 : _GEN_133; 
  assign _GEN_135 = 7'h5 == auto_in_a_bits_source ? _T_499 : _GEN_134; 
  assign _GEN_136 = 7'h6 == auto_in_a_bits_source ? _T_527 : _GEN_135; 
  assign _GEN_137 = 7'h7 == auto_in_a_bits_source ? _T_555 : _GEN_136; 
  assign _GEN_138 = 7'h8 == auto_in_a_bits_source ? _T_583 : _GEN_137; 
  assign _GEN_139 = 7'h9 == auto_in_a_bits_source ? _T_611 : _GEN_138; 
  assign _GEN_140 = 7'ha == auto_in_a_bits_source ? _T_639 : _GEN_139; 
  assign _GEN_141 = 7'hb == auto_in_a_bits_source ? _T_667 : _GEN_140; 
  assign _GEN_142 = 7'hc == auto_in_a_bits_source ? _T_695 : _GEN_141; 
  assign _GEN_143 = 7'hd == auto_in_a_bits_source ? _T_723 : _GEN_142; 
  assign _GEN_144 = 7'he == auto_in_a_bits_source ? _T_751 : _GEN_143; 
  assign _GEN_145 = 7'hf == auto_in_a_bits_source ? _T_779 : _GEN_144; 
  assign _GEN_146 = 7'h10 == auto_in_a_bits_source ? _T_184 : _GEN_145; 
  assign _GEN_147 = 7'h11 == auto_in_a_bits_source ? _T_184 : _GEN_146; 
  assign _GEN_148 = 7'h12 == auto_in_a_bits_source ? _T_184 : _GEN_147; 
  assign _GEN_149 = 7'h13 == auto_in_a_bits_source ? _T_184 : _GEN_148; 
  assign _GEN_150 = 7'h14 == auto_in_a_bits_source ? _T_184 : _GEN_149; 
  assign _GEN_151 = 7'h15 == auto_in_a_bits_source ? _T_184 : _GEN_150; 
  assign _GEN_152 = 7'h16 == auto_in_a_bits_source ? _T_184 : _GEN_151; 
  assign _GEN_153 = 7'h17 == auto_in_a_bits_source ? _T_184 : _GEN_152; 
  assign _GEN_154 = 7'h18 == auto_in_a_bits_source ? _T_184 : _GEN_153; 
  assign _GEN_155 = 7'h19 == auto_in_a_bits_source ? _T_184 : _GEN_154; 
  assign _GEN_156 = 7'h1a == auto_in_a_bits_source ? _T_184 : _GEN_155; 
  assign _GEN_157 = 7'h1b == auto_in_a_bits_source ? _T_184 : _GEN_156; 
  assign _GEN_158 = 7'h1c == auto_in_a_bits_source ? _T_184 : _GEN_157; 
  assign _GEN_159 = 7'h1d == auto_in_a_bits_source ? _T_184 : _GEN_158; 
  assign _GEN_160 = 7'h1e == auto_in_a_bits_source ? _T_184 : _GEN_159; 
  assign _GEN_161 = 7'h1f == auto_in_a_bits_source ? _T_184 : _GEN_160; 
  assign _GEN_162 = 7'h20 == auto_in_a_bits_source ? _T_213 : _GEN_161; 
  assign _GEN_163 = 7'h21 == auto_in_a_bits_source ? _T_213 : _GEN_162; 
  assign _GEN_164 = 7'h22 == auto_in_a_bits_source ? _T_213 : _GEN_163; 
  assign _GEN_165 = 7'h23 == auto_in_a_bits_source ? _T_213 : _GEN_164; 
  assign _GEN_166 = 7'h24 == auto_in_a_bits_source ? _T_213 : _GEN_165; 
  assign _GEN_167 = 7'h25 == auto_in_a_bits_source ? _T_213 : _GEN_166; 
  assign _GEN_168 = 7'h26 == auto_in_a_bits_source ? _T_213 : _GEN_167; 
  assign _GEN_169 = 7'h27 == auto_in_a_bits_source ? _T_213 : _GEN_168; 
  assign _GEN_170 = 7'h28 == auto_in_a_bits_source ? _T_213 : _GEN_169; 
  assign _GEN_171 = 7'h29 == auto_in_a_bits_source ? _T_213 : _GEN_170; 
  assign _GEN_172 = 7'h2a == auto_in_a_bits_source ? _T_213 : _GEN_171; 
  assign _GEN_173 = 7'h2b == auto_in_a_bits_source ? _T_213 : _GEN_172; 
  assign _GEN_174 = 7'h2c == auto_in_a_bits_source ? _T_213 : _GEN_173; 
  assign _GEN_175 = 7'h2d == auto_in_a_bits_source ? _T_213 : _GEN_174; 
  assign _GEN_176 = 7'h2e == auto_in_a_bits_source ? _T_213 : _GEN_175; 
  assign _GEN_177 = 7'h2f == auto_in_a_bits_source ? _T_213 : _GEN_176; 
  assign _GEN_178 = 7'h30 == auto_in_a_bits_source ? _T_242 : _GEN_177; 
  assign _GEN_179 = 7'h31 == auto_in_a_bits_source ? _T_242 : _GEN_178; 
  assign _GEN_180 = 7'h32 == auto_in_a_bits_source ? _T_242 : _GEN_179; 
  assign _GEN_181 = 7'h33 == auto_in_a_bits_source ? _T_242 : _GEN_180; 
  assign _GEN_182 = 7'h34 == auto_in_a_bits_source ? _T_242 : _GEN_181; 
  assign _GEN_183 = 7'h35 == auto_in_a_bits_source ? _T_242 : _GEN_182; 
  assign _GEN_184 = 7'h36 == auto_in_a_bits_source ? _T_242 : _GEN_183; 
  assign _GEN_185 = 7'h37 == auto_in_a_bits_source ? _T_242 : _GEN_184; 
  assign _GEN_186 = 7'h38 == auto_in_a_bits_source ? _T_242 : _GEN_185; 
  assign _GEN_187 = 7'h39 == auto_in_a_bits_source ? _T_242 : _GEN_186; 
  assign _GEN_188 = 7'h3a == auto_in_a_bits_source ? _T_242 : _GEN_187; 
  assign _GEN_189 = 7'h3b == auto_in_a_bits_source ? _T_242 : _GEN_188; 
  assign _GEN_190 = 7'h3c == auto_in_a_bits_source ? _T_242 : _GEN_189; 
  assign _GEN_191 = 7'h3d == auto_in_a_bits_source ? _T_242 : _GEN_190; 
  assign _GEN_192 = 7'h3e == auto_in_a_bits_source ? _T_242 : _GEN_191; 
  assign _GEN_193 = 7'h3f == auto_in_a_bits_source ? _T_242 : _GEN_192; 
  assign _GEN_194 = 7'h40 == auto_in_a_bits_source ? _T_271 : _GEN_193; 
  assign _GEN_195 = 7'h41 == auto_in_a_bits_source ? _T_271 : _GEN_194; 
  assign _GEN_196 = 7'h42 == auto_in_a_bits_source ? _T_271 : _GEN_195; 
  assign _GEN_197 = 7'h43 == auto_in_a_bits_source ? _T_271 : _GEN_196; 
  assign _GEN_198 = 7'h44 == auto_in_a_bits_source ? _T_271 : _GEN_197; 
  assign _GEN_199 = 7'h45 == auto_in_a_bits_source ? _T_271 : _GEN_198; 
  assign _GEN_200 = 7'h46 == auto_in_a_bits_source ? _T_271 : _GEN_199; 
  assign _GEN_201 = 7'h47 == auto_in_a_bits_source ? _T_271 : _GEN_200; 
  assign _GEN_202 = 7'h48 == auto_in_a_bits_source ? _T_271 : _GEN_201; 
  assign _GEN_203 = 7'h49 == auto_in_a_bits_source ? _T_271 : _GEN_202; 
  assign _GEN_204 = 7'h4a == auto_in_a_bits_source ? _T_271 : _GEN_203; 
  assign _GEN_205 = 7'h4b == auto_in_a_bits_source ? _T_271 : _GEN_204; 
  assign _GEN_206 = 7'h4c == auto_in_a_bits_source ? _T_271 : _GEN_205; 
  assign _GEN_207 = 7'h4d == auto_in_a_bits_source ? _T_271 : _GEN_206; 
  assign _GEN_208 = 7'h4e == auto_in_a_bits_source ? _T_271 : _GEN_207; 
  assign _GEN_209 = 7'h4f == auto_in_a_bits_source ? _T_271 : _GEN_208; 
  assign _GEN_210 = 7'h50 == auto_in_a_bits_source ? _T_300 : _GEN_209; 
  assign _GEN_211 = 7'h51 == auto_in_a_bits_source ? _T_300 : _GEN_210; 
  assign _GEN_212 = 7'h52 == auto_in_a_bits_source ? _T_300 : _GEN_211; 
  assign _GEN_213 = 7'h53 == auto_in_a_bits_source ? _T_300 : _GEN_212; 
  assign _GEN_214 = 7'h54 == auto_in_a_bits_source ? _T_300 : _GEN_213; 
  assign _GEN_215 = 7'h55 == auto_in_a_bits_source ? _T_300 : _GEN_214; 
  assign _GEN_216 = 7'h56 == auto_in_a_bits_source ? _T_300 : _GEN_215; 
  assign _GEN_217 = 7'h57 == auto_in_a_bits_source ? _T_300 : _GEN_216; 
  assign _GEN_218 = 7'h58 == auto_in_a_bits_source ? _T_300 : _GEN_217; 
  assign _GEN_219 = 7'h59 == auto_in_a_bits_source ? _T_300 : _GEN_218; 
  assign _GEN_220 = 7'h5a == auto_in_a_bits_source ? _T_300 : _GEN_219; 
  assign _GEN_221 = 7'h5b == auto_in_a_bits_source ? _T_300 : _GEN_220; 
  assign _GEN_222 = 7'h5c == auto_in_a_bits_source ? _T_300 : _GEN_221; 
  assign _GEN_223 = 7'h5d == auto_in_a_bits_source ? _T_300 : _GEN_222; 
  assign _GEN_224 = 7'h5e == auto_in_a_bits_source ? _T_300 : _GEN_223; 
  assign _GEN_225 = 7'h5f == auto_in_a_bits_source ? _T_300 : _GEN_224; 
  assign _GEN_226 = 7'h60 == auto_in_a_bits_source ? _T_329 : _GEN_225; 
  assign _GEN_227 = 7'h61 == auto_in_a_bits_source ? _T_329 : _GEN_226; 
  assign _GEN_228 = 7'h62 == auto_in_a_bits_source ? _T_329 : _GEN_227; 
  assign _GEN_229 = 7'h63 == auto_in_a_bits_source ? _T_329 : _GEN_228; 
  assign _GEN_230 = 7'h64 == auto_in_a_bits_source ? _T_329 : _GEN_229; 
  assign _GEN_231 = 7'h65 == auto_in_a_bits_source ? _T_329 : _GEN_230; 
  assign _GEN_232 = 7'h66 == auto_in_a_bits_source ? _T_329 : _GEN_231; 
  assign _GEN_233 = 7'h67 == auto_in_a_bits_source ? _T_329 : _GEN_232; 
  assign _GEN_234 = 7'h68 == auto_in_a_bits_source ? _T_329 : _GEN_233; 
  assign _GEN_235 = 7'h69 == auto_in_a_bits_source ? _T_329 : _GEN_234; 
  assign _GEN_236 = 7'h6a == auto_in_a_bits_source ? _T_329 : _GEN_235; 
  assign _GEN_237 = 7'h6b == auto_in_a_bits_source ? _T_329 : _GEN_236; 
  assign _GEN_238 = 7'h6c == auto_in_a_bits_source ? _T_329 : _GEN_237; 
  assign _GEN_239 = 7'h6d == auto_in_a_bits_source ? _T_329 : _GEN_238; 
  assign _GEN_240 = 7'h6e == auto_in_a_bits_source ? _T_329 : _GEN_239; 
  assign _GEN_241 = 7'h6f == auto_in_a_bits_source ? _T_329 : _GEN_240; 
  assign _GEN_242 = 7'h70 == auto_in_a_bits_source ? _T_358 : _GEN_241; 
  assign _GEN_243 = 7'h71 == auto_in_a_bits_source ? _T_358 : _GEN_242; 
  assign _GEN_244 = 7'h72 == auto_in_a_bits_source ? _T_358 : _GEN_243; 
  assign _GEN_245 = 7'h73 == auto_in_a_bits_source ? _T_358 : _GEN_244; 
  assign _GEN_246 = 7'h74 == auto_in_a_bits_source ? _T_358 : _GEN_245; 
  assign _GEN_247 = 7'h75 == auto_in_a_bits_source ? _T_358 : _GEN_246; 
  assign _GEN_248 = 7'h76 == auto_in_a_bits_source ? _T_358 : _GEN_247; 
  assign _GEN_249 = 7'h77 == auto_in_a_bits_source ? _T_358 : _GEN_248; 
  assign _GEN_250 = 7'h78 == auto_in_a_bits_source ? _T_358 : _GEN_249; 
  assign _GEN_251 = 7'h79 == auto_in_a_bits_source ? _T_358 : _GEN_250; 
  assign _GEN_252 = 7'h7a == auto_in_a_bits_source ? _T_358 : _GEN_251; 
  assign _GEN_253 = 7'h7b == auto_in_a_bits_source ? _T_358 : _GEN_252; 
  assign _GEN_254 = 7'h7c == auto_in_a_bits_source ? _T_358 : _GEN_253; 
  assign _GEN_255 = 7'h7d == auto_in_a_bits_source ? _T_358 : _GEN_254; 
  assign _GEN_256 = 7'h7e == auto_in_a_bits_source ? _T_358 : _GEN_255; 
  assign _GEN_257 = 7'h7f == auto_in_a_bits_source ? _T_358 : _GEN_256; 
  assign _T_26 = _T_23 == 5'h0; 
  assign _T_67 = _GEN_257 & _T_26; 
  assign _T_68 = _T_67 == 1'h0; 
  assign _T_49_ready = Queue_1_io_enq_ready; 
  assign _T_69 = _T_57 | _T_49_ready; 
  assign _T_50_ready = Queue_io_enq_ready; 
  assign _T_70 = _T_69 & _T_50_ready; 
  assign _T_71 = _T_13 ? _T_70 : _T_49_ready; 
  assign _T_72 = _T_68 & _T_71; 
  assign _T_14 = _T_72 & auto_in_a_valid; 
  assign _T_16 = 23'hff << auto_in_a_bits_size; 
  assign _T_17 = _T_16[7:0]; 
  assign _T_18 = ~ _T_17; 
  assign _T_19 = _T_18[7:3]; 
  assign _T_22 = _T_13 ? _T_19 : 5'h0; 
  assign _T_25 = _T_23 - 5'h1; 
  assign _T_27 = _T_23 == 5'h1; 
  assign _T_28 = _T_22 == 5'h0; 
  assign _T_29 = _T_27 | _T_28; 
  assign _T_43 = {auto_in_a_bits_size, 7'h0}; 
  assign _GEN_284 = {{4'd0}, auto_in_a_bits_source}; 
  assign _T_45 = auto_out_ruser[6:0]; 
  assign _T_46 = auto_out_ruser[10:7]; 
  assign _T_47 = auto_out_buser[6:0]; 
  assign _T_48 = auto_out_buser[10:7]; 
  assign _T_52_bits_wen = Queue_1_io_deq_bits_wen; 
  assign _T_53 = _T_52_bits_wen == 1'h0; 
  assign _T_52_valid = Queue_1_io_deq_valid; 
  assign _T_59 = _T_29 == 1'h0; 
  assign _GEN_3 = 7'h1 == auto_in_a_bits_source ? 5'h8 : 5'h7; 
  assign _GEN_4 = 7'h2 == auto_in_a_bits_source ? 5'h9 : _GEN_3; 
  assign _GEN_5 = 7'h3 == auto_in_a_bits_source ? 5'ha : _GEN_4; 
  assign _GEN_6 = 7'h4 == auto_in_a_bits_source ? 5'hb : _GEN_5; 
  assign _GEN_7 = 7'h5 == auto_in_a_bits_source ? 5'hc : _GEN_6; 
  assign _GEN_8 = 7'h6 == auto_in_a_bits_source ? 5'hd : _GEN_7; 
  assign _GEN_9 = 7'h7 == auto_in_a_bits_source ? 5'he : _GEN_8; 
  assign _GEN_10 = 7'h8 == auto_in_a_bits_source ? 5'hf : _GEN_9; 
  assign _GEN_11 = 7'h9 == auto_in_a_bits_source ? 5'h10 : _GEN_10; 
  assign _GEN_12 = 7'ha == auto_in_a_bits_source ? 5'h11 : _GEN_11; 
  assign _GEN_13 = 7'hb == auto_in_a_bits_source ? 5'h12 : _GEN_12; 
  assign _GEN_14 = 7'hc == auto_in_a_bits_source ? 5'h13 : _GEN_13; 
  assign _GEN_15 = 7'hd == auto_in_a_bits_source ? 5'h14 : _GEN_14; 
  assign _GEN_16 = 7'he == auto_in_a_bits_source ? 5'h15 : _GEN_15; 
  assign _GEN_17 = 7'hf == auto_in_a_bits_source ? 5'h16 : _GEN_16; 
  assign _GEN_18 = 7'h10 == auto_in_a_bits_source ? 5'h0 : _GEN_17; 
  assign _GEN_19 = 7'h11 == auto_in_a_bits_source ? 5'h0 : _GEN_18; 
  assign _GEN_20 = 7'h12 == auto_in_a_bits_source ? 5'h0 : _GEN_19; 
  assign _GEN_21 = 7'h13 == auto_in_a_bits_source ? 5'h0 : _GEN_20; 
  assign _GEN_22 = 7'h14 == auto_in_a_bits_source ? 5'h0 : _GEN_21; 
  assign _GEN_23 = 7'h15 == auto_in_a_bits_source ? 5'h0 : _GEN_22; 
  assign _GEN_24 = 7'h16 == auto_in_a_bits_source ? 5'h0 : _GEN_23; 
  assign _GEN_25 = 7'h17 == auto_in_a_bits_source ? 5'h0 : _GEN_24; 
  assign _GEN_26 = 7'h18 == auto_in_a_bits_source ? 5'h0 : _GEN_25; 
  assign _GEN_27 = 7'h19 == auto_in_a_bits_source ? 5'h0 : _GEN_26; 
  assign _GEN_28 = 7'h1a == auto_in_a_bits_source ? 5'h0 : _GEN_27; 
  assign _GEN_29 = 7'h1b == auto_in_a_bits_source ? 5'h0 : _GEN_28; 
  assign _GEN_30 = 7'h1c == auto_in_a_bits_source ? 5'h0 : _GEN_29; 
  assign _GEN_31 = 7'h1d == auto_in_a_bits_source ? 5'h0 : _GEN_30; 
  assign _GEN_32 = 7'h1e == auto_in_a_bits_source ? 5'h0 : _GEN_31; 
  assign _GEN_33 = 7'h1f == auto_in_a_bits_source ? 5'h0 : _GEN_32; 
  assign _GEN_34 = 7'h20 == auto_in_a_bits_source ? 5'h1 : _GEN_33; 
  assign _GEN_35 = 7'h21 == auto_in_a_bits_source ? 5'h1 : _GEN_34; 
  assign _GEN_36 = 7'h22 == auto_in_a_bits_source ? 5'h1 : _GEN_35; 
  assign _GEN_37 = 7'h23 == auto_in_a_bits_source ? 5'h1 : _GEN_36; 
  assign _GEN_38 = 7'h24 == auto_in_a_bits_source ? 5'h1 : _GEN_37; 
  assign _GEN_39 = 7'h25 == auto_in_a_bits_source ? 5'h1 : _GEN_38; 
  assign _GEN_40 = 7'h26 == auto_in_a_bits_source ? 5'h1 : _GEN_39; 
  assign _GEN_41 = 7'h27 == auto_in_a_bits_source ? 5'h1 : _GEN_40; 
  assign _GEN_42 = 7'h28 == auto_in_a_bits_source ? 5'h1 : _GEN_41; 
  assign _GEN_43 = 7'h29 == auto_in_a_bits_source ? 5'h1 : _GEN_42; 
  assign _GEN_44 = 7'h2a == auto_in_a_bits_source ? 5'h1 : _GEN_43; 
  assign _GEN_45 = 7'h2b == auto_in_a_bits_source ? 5'h1 : _GEN_44; 
  assign _GEN_46 = 7'h2c == auto_in_a_bits_source ? 5'h1 : _GEN_45; 
  assign _GEN_47 = 7'h2d == auto_in_a_bits_source ? 5'h1 : _GEN_46; 
  assign _GEN_48 = 7'h2e == auto_in_a_bits_source ? 5'h1 : _GEN_47; 
  assign _GEN_49 = 7'h2f == auto_in_a_bits_source ? 5'h1 : _GEN_48; 
  assign _GEN_50 = 7'h30 == auto_in_a_bits_source ? 5'h2 : _GEN_49; 
  assign _GEN_51 = 7'h31 == auto_in_a_bits_source ? 5'h2 : _GEN_50; 
  assign _GEN_52 = 7'h32 == auto_in_a_bits_source ? 5'h2 : _GEN_51; 
  assign _GEN_53 = 7'h33 == auto_in_a_bits_source ? 5'h2 : _GEN_52; 
  assign _GEN_54 = 7'h34 == auto_in_a_bits_source ? 5'h2 : _GEN_53; 
  assign _GEN_55 = 7'h35 == auto_in_a_bits_source ? 5'h2 : _GEN_54; 
  assign _GEN_56 = 7'h36 == auto_in_a_bits_source ? 5'h2 : _GEN_55; 
  assign _GEN_57 = 7'h37 == auto_in_a_bits_source ? 5'h2 : _GEN_56; 
  assign _GEN_58 = 7'h38 == auto_in_a_bits_source ? 5'h2 : _GEN_57; 
  assign _GEN_59 = 7'h39 == auto_in_a_bits_source ? 5'h2 : _GEN_58; 
  assign _GEN_60 = 7'h3a == auto_in_a_bits_source ? 5'h2 : _GEN_59; 
  assign _GEN_61 = 7'h3b == auto_in_a_bits_source ? 5'h2 : _GEN_60; 
  assign _GEN_62 = 7'h3c == auto_in_a_bits_source ? 5'h2 : _GEN_61; 
  assign _GEN_63 = 7'h3d == auto_in_a_bits_source ? 5'h2 : _GEN_62; 
  assign _GEN_64 = 7'h3e == auto_in_a_bits_source ? 5'h2 : _GEN_63; 
  assign _GEN_65 = 7'h3f == auto_in_a_bits_source ? 5'h2 : _GEN_64; 
  assign _GEN_66 = 7'h40 == auto_in_a_bits_source ? 5'h3 : _GEN_65; 
  assign _GEN_67 = 7'h41 == auto_in_a_bits_source ? 5'h3 : _GEN_66; 
  assign _GEN_68 = 7'h42 == auto_in_a_bits_source ? 5'h3 : _GEN_67; 
  assign _GEN_69 = 7'h43 == auto_in_a_bits_source ? 5'h3 : _GEN_68; 
  assign _GEN_70 = 7'h44 == auto_in_a_bits_source ? 5'h3 : _GEN_69; 
  assign _GEN_71 = 7'h45 == auto_in_a_bits_source ? 5'h3 : _GEN_70; 
  assign _GEN_72 = 7'h46 == auto_in_a_bits_source ? 5'h3 : _GEN_71; 
  assign _GEN_73 = 7'h47 == auto_in_a_bits_source ? 5'h3 : _GEN_72; 
  assign _GEN_74 = 7'h48 == auto_in_a_bits_source ? 5'h3 : _GEN_73; 
  assign _GEN_75 = 7'h49 == auto_in_a_bits_source ? 5'h3 : _GEN_74; 
  assign _GEN_76 = 7'h4a == auto_in_a_bits_source ? 5'h3 : _GEN_75; 
  assign _GEN_77 = 7'h4b == auto_in_a_bits_source ? 5'h3 : _GEN_76; 
  assign _GEN_78 = 7'h4c == auto_in_a_bits_source ? 5'h3 : _GEN_77; 
  assign _GEN_79 = 7'h4d == auto_in_a_bits_source ? 5'h3 : _GEN_78; 
  assign _GEN_80 = 7'h4e == auto_in_a_bits_source ? 5'h3 : _GEN_79; 
  assign _GEN_81 = 7'h4f == auto_in_a_bits_source ? 5'h3 : _GEN_80; 
  assign _GEN_82 = 7'h50 == auto_in_a_bits_source ? 5'h4 : _GEN_81; 
  assign _GEN_83 = 7'h51 == auto_in_a_bits_source ? 5'h4 : _GEN_82; 
  assign _GEN_84 = 7'h52 == auto_in_a_bits_source ? 5'h4 : _GEN_83; 
  assign _GEN_85 = 7'h53 == auto_in_a_bits_source ? 5'h4 : _GEN_84; 
  assign _GEN_86 = 7'h54 == auto_in_a_bits_source ? 5'h4 : _GEN_85; 
  assign _GEN_87 = 7'h55 == auto_in_a_bits_source ? 5'h4 : _GEN_86; 
  assign _GEN_88 = 7'h56 == auto_in_a_bits_source ? 5'h4 : _GEN_87; 
  assign _GEN_89 = 7'h57 == auto_in_a_bits_source ? 5'h4 : _GEN_88; 
  assign _GEN_90 = 7'h58 == auto_in_a_bits_source ? 5'h4 : _GEN_89; 
  assign _GEN_91 = 7'h59 == auto_in_a_bits_source ? 5'h4 : _GEN_90; 
  assign _GEN_92 = 7'h5a == auto_in_a_bits_source ? 5'h4 : _GEN_91; 
  assign _GEN_93 = 7'h5b == auto_in_a_bits_source ? 5'h4 : _GEN_92; 
  assign _GEN_94 = 7'h5c == auto_in_a_bits_source ? 5'h4 : _GEN_93; 
  assign _GEN_95 = 7'h5d == auto_in_a_bits_source ? 5'h4 : _GEN_94; 
  assign _GEN_96 = 7'h5e == auto_in_a_bits_source ? 5'h4 : _GEN_95; 
  assign _GEN_97 = 7'h5f == auto_in_a_bits_source ? 5'h4 : _GEN_96; 
  assign _GEN_98 = 7'h60 == auto_in_a_bits_source ? 5'h5 : _GEN_97; 
  assign _GEN_99 = 7'h61 == auto_in_a_bits_source ? 5'h5 : _GEN_98; 
  assign _GEN_100 = 7'h62 == auto_in_a_bits_source ? 5'h5 : _GEN_99; 
  assign _GEN_101 = 7'h63 == auto_in_a_bits_source ? 5'h5 : _GEN_100; 
  assign _GEN_102 = 7'h64 == auto_in_a_bits_source ? 5'h5 : _GEN_101; 
  assign _GEN_103 = 7'h65 == auto_in_a_bits_source ? 5'h5 : _GEN_102; 
  assign _GEN_104 = 7'h66 == auto_in_a_bits_source ? 5'h5 : _GEN_103; 
  assign _GEN_105 = 7'h67 == auto_in_a_bits_source ? 5'h5 : _GEN_104; 
  assign _GEN_106 = 7'h68 == auto_in_a_bits_source ? 5'h5 : _GEN_105; 
  assign _GEN_107 = 7'h69 == auto_in_a_bits_source ? 5'h5 : _GEN_106; 
  assign _GEN_108 = 7'h6a == auto_in_a_bits_source ? 5'h5 : _GEN_107; 
  assign _GEN_109 = 7'h6b == auto_in_a_bits_source ? 5'h5 : _GEN_108; 
  assign _GEN_110 = 7'h6c == auto_in_a_bits_source ? 5'h5 : _GEN_109; 
  assign _GEN_111 = 7'h6d == auto_in_a_bits_source ? 5'h5 : _GEN_110; 
  assign _GEN_112 = 7'h6e == auto_in_a_bits_source ? 5'h5 : _GEN_111; 
  assign _GEN_113 = 7'h6f == auto_in_a_bits_source ? 5'h5 : _GEN_112; 
  assign _GEN_114 = 7'h70 == auto_in_a_bits_source ? 5'h6 : _GEN_113; 
  assign _GEN_115 = 7'h71 == auto_in_a_bits_source ? 5'h6 : _GEN_114; 
  assign _GEN_116 = 7'h72 == auto_in_a_bits_source ? 5'h6 : _GEN_115; 
  assign _GEN_117 = 7'h73 == auto_in_a_bits_source ? 5'h6 : _GEN_116; 
  assign _GEN_118 = 7'h74 == auto_in_a_bits_source ? 5'h6 : _GEN_117; 
  assign _GEN_119 = 7'h75 == auto_in_a_bits_source ? 5'h6 : _GEN_118; 
  assign _GEN_120 = 7'h76 == auto_in_a_bits_source ? 5'h6 : _GEN_119; 
  assign _GEN_121 = 7'h77 == auto_in_a_bits_source ? 5'h6 : _GEN_120; 
  assign _GEN_122 = 7'h78 == auto_in_a_bits_source ? 5'h6 : _GEN_121; 
  assign _GEN_123 = 7'h79 == auto_in_a_bits_source ? 5'h6 : _GEN_122; 
  assign _GEN_124 = 7'h7a == auto_in_a_bits_source ? 5'h6 : _GEN_123; 
  assign _GEN_125 = 7'h7b == auto_in_a_bits_source ? 5'h6 : _GEN_124; 
  assign _GEN_126 = 7'h7c == auto_in_a_bits_source ? 5'h6 : _GEN_125; 
  assign _GEN_127 = 7'h7d == auto_in_a_bits_source ? 5'h6 : _GEN_126; 
  assign _GEN_128 = 7'h7e == auto_in_a_bits_source ? 5'h6 : _GEN_127; 
  assign _GEN_129 = 7'h7f == auto_in_a_bits_source ? 5'h6 : _GEN_128; 
  assign _T_61 = 26'h7ff << auto_in_a_bits_size; 
  assign _T_62 = _T_61[10:0]; 
  assign _T_63 = ~ _T_62; 
  assign _T_65 = auto_in_a_bits_size >= 4'h3; 
  assign _T_66 = _T_65 ? 4'h3 : auto_in_a_bits_size; 
  assign _T_74 = _T_68 & auto_in_a_valid; 
  assign _T_75 = _T_57 == 1'h0; 
  assign _T_76 = _T_75 & _T_50_ready; 
  assign _T_77 = _T_13 ? _T_76 : 1'h1; 
  assign _T_78 = _T_74 & _T_77; 
  assign _T_81 = _T_74 & _T_13; 
  assign _T_85 = auto_in_d_ready & auto_out_rvalid; 
  assign _T_86 = auto_out_rlast == 1'h0; 
  assign _T_87 = auto_out_rvalid | _T_84; 
  assign _T_88 = _T_87 == 1'h0; 
  assign _T_90 = _T_87 ? auto_out_rvalid : auto_out_bvalid; 
  assign _T_93 = auto_out_rresp == 2'h3; 
  assign _GEN_260 = _T_91 ? _T_93 : _T_94; 
  assign _T_96 = auto_out_rresp != 2'h0; 
  assign _T_97 = auto_out_bresp != 2'h0; 
  assign _T_98 = _T_96 | _GEN_260; 
  assign _T_103 = 32'h1 << _GEN_129; 
  assign _T_104 = _T_103[22:0]; 
  assign _T_105 = _T_104[0]; 
  assign _T_106 = _T_104[1]; 
  assign _T_107 = _T_104[2]; 
  assign _T_108 = _T_104[3]; 
  assign _T_109 = _T_104[4]; 
  assign _T_110 = _T_104[5]; 
  assign _T_111 = _T_104[6]; 
  assign _T_112 = _T_104[7]; 
  assign _T_113 = _T_104[8]; 
  assign _T_114 = _T_104[9]; 
  assign _T_115 = _T_104[10]; 
  assign _T_116 = _T_104[11]; 
  assign _T_117 = _T_104[12]; 
  assign _T_118 = _T_104[13]; 
  assign _T_119 = _T_104[14]; 
  assign _T_120 = _T_104[15]; 
  assign _T_121 = _T_104[16]; 
  assign _T_122 = _T_104[17]; 
  assign _T_123 = _T_104[18]; 
  assign _T_124 = _T_104[19]; 
  assign _T_125 = _T_104[20]; 
  assign _T_126 = _T_104[21]; 
  assign _T_127 = _T_104[22]; 
  assign _T_128 = _T_87 ? auto_out_rid : auto_out_bid; 
  assign _T_130 = 32'h1 << _T_128; 
  assign _T_131 = _T_130[22:0]; 
  assign _T_132 = _T_131[0]; 
  assign _T_133 = _T_131[1]; 
  assign _T_134 = _T_131[2]; 
  assign _T_135 = _T_131[3]; 
  assign _T_136 = _T_131[4]; 
  assign _T_137 = _T_131[5]; 
  assign _T_138 = _T_131[6]; 
  assign _T_139 = _T_131[7]; 
  assign _T_140 = _T_131[8]; 
  assign _T_141 = _T_131[9]; 
  assign _T_142 = _T_131[10]; 
  assign _T_143 = _T_131[11]; 
  assign _T_144 = _T_131[12]; 
  assign _T_145 = _T_131[13]; 
  assign _T_146 = _T_131[14]; 
  assign _T_147 = _T_131[15]; 
  assign _T_148 = _T_131[16]; 
  assign _T_149 = _T_131[17]; 
  assign _T_150 = _T_131[18]; 
  assign _T_151 = _T_131[19]; 
  assign _T_152 = _T_131[20]; 
  assign _T_153 = _T_131[21]; 
  assign _T_154 = _T_131[22]; 
  assign _T_155 = _T_87 ? auto_out_rlast : 1'h1; 
  assign _T_159 = _T_49_ready & _T_78; 
  assign _T_160 = _T_105 & _T_159; 
  assign _T_161 = _T_132 & _T_155; 
  assign _T_162 = auto_in_d_ready & _T_90; 
  assign _T_163 = _T_161 & _T_162; 
  assign _GEN_285 = {{4'd0}, _T_160}; 
  assign _T_165 = _T_156 + _GEN_285; 
  assign _GEN_286 = {{4'd0}, _T_163}; 
  assign _T_167 = _T_165 - _GEN_286; 
  assign _T_168 = _T_163 == 1'h0; 
  assign _T_169 = _T_156 != 5'h0; 
  assign _T_170 = _T_168 | _T_169; 
  assign _T_172 = _T_170 | reset; 
  assign _T_173 = _T_172 == 1'h0; 
  assign _T_174 = _T_160 == 1'h0; 
  assign _T_175 = _T_156 != 5'h10; 
  assign _T_176 = _T_174 | _T_175; 
  assign _T_178 = _T_176 | reset; 
  assign _T_179 = _T_178 == 1'h0; 
  assign _T_189 = _T_106 & _T_159; 
  assign _T_190 = _T_133 & _T_155; 
  assign _T_192 = _T_190 & _T_162; 
  assign _GEN_287 = {{4'd0}, _T_189}; 
  assign _T_194 = _T_185 + _GEN_287; 
  assign _GEN_288 = {{4'd0}, _T_192}; 
  assign _T_196 = _T_194 - _GEN_288; 
  assign _T_197 = _T_192 == 1'h0; 
  assign _T_198 = _T_185 != 5'h0; 
  assign _T_199 = _T_197 | _T_198; 
  assign _T_201 = _T_199 | reset; 
  assign _T_202 = _T_201 == 1'h0; 
  assign _T_203 = _T_189 == 1'h0; 
  assign _T_204 = _T_185 != 5'h10; 
  assign _T_205 = _T_203 | _T_204; 
  assign _T_207 = _T_205 | reset; 
  assign _T_208 = _T_207 == 1'h0; 
  assign _T_218 = _T_107 & _T_159; 
  assign _T_219 = _T_134 & _T_155; 
  assign _T_221 = _T_219 & _T_162; 
  assign _GEN_289 = {{4'd0}, _T_218}; 
  assign _T_223 = _T_214 + _GEN_289; 
  assign _GEN_290 = {{4'd0}, _T_221}; 
  assign _T_225 = _T_223 - _GEN_290; 
  assign _T_226 = _T_221 == 1'h0; 
  assign _T_227 = _T_214 != 5'h0; 
  assign _T_228 = _T_226 | _T_227; 
  assign _T_230 = _T_228 | reset; 
  assign _T_231 = _T_230 == 1'h0; 
  assign _T_232 = _T_218 == 1'h0; 
  assign _T_233 = _T_214 != 5'h10; 
  assign _T_234 = _T_232 | _T_233; 
  assign _T_236 = _T_234 | reset; 
  assign _T_237 = _T_236 == 1'h0; 
  assign _T_247 = _T_108 & _T_159; 
  assign _T_248 = _T_135 & _T_155; 
  assign _T_250 = _T_248 & _T_162; 
  assign _GEN_291 = {{4'd0}, _T_247}; 
  assign _T_252 = _T_243 + _GEN_291; 
  assign _GEN_292 = {{4'd0}, _T_250}; 
  assign _T_254 = _T_252 - _GEN_292; 
  assign _T_255 = _T_250 == 1'h0; 
  assign _T_256 = _T_243 != 5'h0; 
  assign _T_257 = _T_255 | _T_256; 
  assign _T_259 = _T_257 | reset; 
  assign _T_260 = _T_259 == 1'h0; 
  assign _T_261 = _T_247 == 1'h0; 
  assign _T_262 = _T_243 != 5'h10; 
  assign _T_263 = _T_261 | _T_262; 
  assign _T_265 = _T_263 | reset; 
  assign _T_266 = _T_265 == 1'h0; 
  assign _T_276 = _T_109 & _T_159; 
  assign _T_277 = _T_136 & _T_155; 
  assign _T_279 = _T_277 & _T_162; 
  assign _GEN_293 = {{4'd0}, _T_276}; 
  assign _T_281 = _T_272 + _GEN_293; 
  assign _GEN_294 = {{4'd0}, _T_279}; 
  assign _T_283 = _T_281 - _GEN_294; 
  assign _T_284 = _T_279 == 1'h0; 
  assign _T_285 = _T_272 != 5'h0; 
  assign _T_286 = _T_284 | _T_285; 
  assign _T_288 = _T_286 | reset; 
  assign _T_289 = _T_288 == 1'h0; 
  assign _T_290 = _T_276 == 1'h0; 
  assign _T_291 = _T_272 != 5'h10; 
  assign _T_292 = _T_290 | _T_291; 
  assign _T_294 = _T_292 | reset; 
  assign _T_295 = _T_294 == 1'h0; 
  assign _T_305 = _T_110 & _T_159; 
  assign _T_306 = _T_137 & _T_155; 
  assign _T_308 = _T_306 & _T_162; 
  assign _GEN_295 = {{4'd0}, _T_305}; 
  assign _T_310 = _T_301 + _GEN_295; 
  assign _GEN_296 = {{4'd0}, _T_308}; 
  assign _T_312 = _T_310 - _GEN_296; 
  assign _T_313 = _T_308 == 1'h0; 
  assign _T_314 = _T_301 != 5'h0; 
  assign _T_315 = _T_313 | _T_314; 
  assign _T_317 = _T_315 | reset; 
  assign _T_318 = _T_317 == 1'h0; 
  assign _T_319 = _T_305 == 1'h0; 
  assign _T_320 = _T_301 != 5'h10; 
  assign _T_321 = _T_319 | _T_320; 
  assign _T_323 = _T_321 | reset; 
  assign _T_324 = _T_323 == 1'h0; 
  assign _T_334 = _T_111 & _T_159; 
  assign _T_335 = _T_138 & _T_155; 
  assign _T_337 = _T_335 & _T_162; 
  assign _GEN_297 = {{4'd0}, _T_334}; 
  assign _T_339 = _T_330 + _GEN_297; 
  assign _GEN_298 = {{4'd0}, _T_337}; 
  assign _T_341 = _T_339 - _GEN_298; 
  assign _T_342 = _T_337 == 1'h0; 
  assign _T_343 = _T_330 != 5'h0; 
  assign _T_344 = _T_342 | _T_343; 
  assign _T_346 = _T_344 | reset; 
  assign _T_347 = _T_346 == 1'h0; 
  assign _T_348 = _T_334 == 1'h0; 
  assign _T_349 = _T_330 != 5'h10; 
  assign _T_350 = _T_348 | _T_349; 
  assign _T_352 = _T_350 | reset; 
  assign _T_353 = _T_352 == 1'h0; 
  assign _T_363 = _T_112 & _T_159; 
  assign _T_364 = _T_139 & _T_155; 
  assign _T_366 = _T_364 & _T_162; 
  assign _T_368 = _T_359 + _T_363; 
  assign _T_370 = _T_368 - _T_366; 
  assign _T_371 = _T_366 == 1'h0; 
  assign _T_373 = _T_371 | _T_359; 
  assign _T_375 = _T_373 | reset; 
  assign _T_376 = _T_375 == 1'h0; 
  assign _T_377 = _T_363 == 1'h0; 
  assign _T_378 = _T_359 != 1'h1; 
  assign _T_379 = _T_377 | _T_378; 
  assign _T_381 = _T_379 | reset; 
  assign _T_382 = _T_381 == 1'h0; 
  assign _T_391 = _T_113 & _T_159; 
  assign _T_392 = _T_140 & _T_155; 
  assign _T_394 = _T_392 & _T_162; 
  assign _T_396 = _T_387 + _T_391; 
  assign _T_398 = _T_396 - _T_394; 
  assign _T_399 = _T_394 == 1'h0; 
  assign _T_401 = _T_399 | _T_387; 
  assign _T_403 = _T_401 | reset; 
  assign _T_404 = _T_403 == 1'h0; 
  assign _T_405 = _T_391 == 1'h0; 
  assign _T_406 = _T_387 != 1'h1; 
  assign _T_407 = _T_405 | _T_406; 
  assign _T_409 = _T_407 | reset; 
  assign _T_410 = _T_409 == 1'h0; 
  assign _T_419 = _T_114 & _T_159; 
  assign _T_420 = _T_141 & _T_155; 
  assign _T_422 = _T_420 & _T_162; 
  assign _T_424 = _T_415 + _T_419; 
  assign _T_426 = _T_424 - _T_422; 
  assign _T_427 = _T_422 == 1'h0; 
  assign _T_429 = _T_427 | _T_415; 
  assign _T_431 = _T_429 | reset; 
  assign _T_432 = _T_431 == 1'h0; 
  assign _T_433 = _T_419 == 1'h0; 
  assign _T_434 = _T_415 != 1'h1; 
  assign _T_435 = _T_433 | _T_434; 
  assign _T_437 = _T_435 | reset; 
  assign _T_438 = _T_437 == 1'h0; 
  assign _T_447 = _T_115 & _T_159; 
  assign _T_448 = _T_142 & _T_155; 
  assign _T_450 = _T_448 & _T_162; 
  assign _T_452 = _T_443 + _T_447; 
  assign _T_454 = _T_452 - _T_450; 
  assign _T_455 = _T_450 == 1'h0; 
  assign _T_457 = _T_455 | _T_443; 
  assign _T_459 = _T_457 | reset; 
  assign _T_460 = _T_459 == 1'h0; 
  assign _T_461 = _T_447 == 1'h0; 
  assign _T_462 = _T_443 != 1'h1; 
  assign _T_463 = _T_461 | _T_462; 
  assign _T_465 = _T_463 | reset; 
  assign _T_466 = _T_465 == 1'h0; 
  assign _T_475 = _T_116 & _T_159; 
  assign _T_476 = _T_143 & _T_155; 
  assign _T_478 = _T_476 & _T_162; 
  assign _T_480 = _T_471 + _T_475; 
  assign _T_482 = _T_480 - _T_478; 
  assign _T_483 = _T_478 == 1'h0; 
  assign _T_485 = _T_483 | _T_471; 
  assign _T_487 = _T_485 | reset; 
  assign _T_488 = _T_487 == 1'h0; 
  assign _T_489 = _T_475 == 1'h0; 
  assign _T_490 = _T_471 != 1'h1; 
  assign _T_491 = _T_489 | _T_490; 
  assign _T_493 = _T_491 | reset; 
  assign _T_494 = _T_493 == 1'h0; 
  assign _T_503 = _T_117 & _T_159; 
  assign _T_504 = _T_144 & _T_155; 
  assign _T_506 = _T_504 & _T_162; 
  assign _T_508 = _T_499 + _T_503; 
  assign _T_510 = _T_508 - _T_506; 
  assign _T_511 = _T_506 == 1'h0; 
  assign _T_513 = _T_511 | _T_499; 
  assign _T_515 = _T_513 | reset; 
  assign _T_516 = _T_515 == 1'h0; 
  assign _T_517 = _T_503 == 1'h0; 
  assign _T_518 = _T_499 != 1'h1; 
  assign _T_519 = _T_517 | _T_518; 
  assign _T_521 = _T_519 | reset; 
  assign _T_522 = _T_521 == 1'h0; 
  assign _T_531 = _T_118 & _T_159; 
  assign _T_532 = _T_145 & _T_155; 
  assign _T_534 = _T_532 & _T_162; 
  assign _T_536 = _T_527 + _T_531; 
  assign _T_538 = _T_536 - _T_534; 
  assign _T_539 = _T_534 == 1'h0; 
  assign _T_541 = _T_539 | _T_527; 
  assign _T_543 = _T_541 | reset; 
  assign _T_544 = _T_543 == 1'h0; 
  assign _T_545 = _T_531 == 1'h0; 
  assign _T_546 = _T_527 != 1'h1; 
  assign _T_547 = _T_545 | _T_546; 
  assign _T_549 = _T_547 | reset; 
  assign _T_550 = _T_549 == 1'h0; 
  assign _T_559 = _T_119 & _T_159; 
  assign _T_560 = _T_146 & _T_155; 
  assign _T_562 = _T_560 & _T_162; 
  assign _T_564 = _T_555 + _T_559; 
  assign _T_566 = _T_564 - _T_562; 
  assign _T_567 = _T_562 == 1'h0; 
  assign _T_569 = _T_567 | _T_555; 
  assign _T_571 = _T_569 | reset; 
  assign _T_572 = _T_571 == 1'h0; 
  assign _T_573 = _T_559 == 1'h0; 
  assign _T_574 = _T_555 != 1'h1; 
  assign _T_575 = _T_573 | _T_574; 
  assign _T_577 = _T_575 | reset; 
  assign _T_578 = _T_577 == 1'h0; 
  assign _T_587 = _T_120 & _T_159; 
  assign _T_588 = _T_147 & _T_155; 
  assign _T_590 = _T_588 & _T_162; 
  assign _T_592 = _T_583 + _T_587; 
  assign _T_594 = _T_592 - _T_590; 
  assign _T_595 = _T_590 == 1'h0; 
  assign _T_597 = _T_595 | _T_583; 
  assign _T_599 = _T_597 | reset; 
  assign _T_600 = _T_599 == 1'h0; 
  assign _T_601 = _T_587 == 1'h0; 
  assign _T_602 = _T_583 != 1'h1; 
  assign _T_603 = _T_601 | _T_602; 
  assign _T_605 = _T_603 | reset; 
  assign _T_606 = _T_605 == 1'h0; 
  assign _T_615 = _T_121 & _T_159; 
  assign _T_616 = _T_148 & _T_155; 
  assign _T_618 = _T_616 & _T_162; 
  assign _T_620 = _T_611 + _T_615; 
  assign _T_622 = _T_620 - _T_618; 
  assign _T_623 = _T_618 == 1'h0; 
  assign _T_625 = _T_623 | _T_611; 
  assign _T_627 = _T_625 | reset; 
  assign _T_628 = _T_627 == 1'h0; 
  assign _T_629 = _T_615 == 1'h0; 
  assign _T_630 = _T_611 != 1'h1; 
  assign _T_631 = _T_629 | _T_630; 
  assign _T_633 = _T_631 | reset; 
  assign _T_634 = _T_633 == 1'h0; 
  assign _T_643 = _T_122 & _T_159; 
  assign _T_644 = _T_149 & _T_155; 
  assign _T_646 = _T_644 & _T_162; 
  assign _T_648 = _T_639 + _T_643; 
  assign _T_650 = _T_648 - _T_646; 
  assign _T_651 = _T_646 == 1'h0; 
  assign _T_653 = _T_651 | _T_639; 
  assign _T_655 = _T_653 | reset; 
  assign _T_656 = _T_655 == 1'h0; 
  assign _T_657 = _T_643 == 1'h0; 
  assign _T_658 = _T_639 != 1'h1; 
  assign _T_659 = _T_657 | _T_658; 
  assign _T_661 = _T_659 | reset; 
  assign _T_662 = _T_661 == 1'h0; 
  assign _T_671 = _T_123 & _T_159; 
  assign _T_672 = _T_150 & _T_155; 
  assign _T_674 = _T_672 & _T_162; 
  assign _T_676 = _T_667 + _T_671; 
  assign _T_678 = _T_676 - _T_674; 
  assign _T_679 = _T_674 == 1'h0; 
  assign _T_681 = _T_679 | _T_667; 
  assign _T_683 = _T_681 | reset; 
  assign _T_684 = _T_683 == 1'h0; 
  assign _T_685 = _T_671 == 1'h0; 
  assign _T_686 = _T_667 != 1'h1; 
  assign _T_687 = _T_685 | _T_686; 
  assign _T_689 = _T_687 | reset; 
  assign _T_690 = _T_689 == 1'h0; 
  assign _T_699 = _T_124 & _T_159; 
  assign _T_700 = _T_151 & _T_155; 
  assign _T_702 = _T_700 & _T_162; 
  assign _T_704 = _T_695 + _T_699; 
  assign _T_706 = _T_704 - _T_702; 
  assign _T_707 = _T_702 == 1'h0; 
  assign _T_709 = _T_707 | _T_695; 
  assign _T_711 = _T_709 | reset; 
  assign _T_712 = _T_711 == 1'h0; 
  assign _T_713 = _T_699 == 1'h0; 
  assign _T_714 = _T_695 != 1'h1; 
  assign _T_715 = _T_713 | _T_714; 
  assign _T_717 = _T_715 | reset; 
  assign _T_718 = _T_717 == 1'h0; 
  assign _T_727 = _T_125 & _T_159; 
  assign _T_728 = _T_152 & _T_155; 
  assign _T_730 = _T_728 & _T_162; 
  assign _T_732 = _T_723 + _T_727; 
  assign _T_734 = _T_732 - _T_730; 
  assign _T_735 = _T_730 == 1'h0; 
  assign _T_737 = _T_735 | _T_723; 
  assign _T_739 = _T_737 | reset; 
  assign _T_740 = _T_739 == 1'h0; 
  assign _T_741 = _T_727 == 1'h0; 
  assign _T_742 = _T_723 != 1'h1; 
  assign _T_743 = _T_741 | _T_742; 
  assign _T_745 = _T_743 | reset; 
  assign _T_746 = _T_745 == 1'h0; 
  assign _T_755 = _T_126 & _T_159; 
  assign _T_756 = _T_153 & _T_155; 
  assign _T_758 = _T_756 & _T_162; 
  assign _T_760 = _T_751 + _T_755; 
  assign _T_762 = _T_760 - _T_758; 
  assign _T_763 = _T_758 == 1'h0; 
  assign _T_765 = _T_763 | _T_751; 
  assign _T_767 = _T_765 | reset; 
  assign _T_768 = _T_767 == 1'h0; 
  assign _T_769 = _T_755 == 1'h0; 
  assign _T_770 = _T_751 != 1'h1; 
  assign _T_771 = _T_769 | _T_770; 
  assign _T_773 = _T_771 | reset; 
  assign _T_774 = _T_773 == 1'h0; 
  assign _T_783 = _T_127 & _T_159; 
  assign _T_784 = _T_154 & _T_155; 
  assign _T_786 = _T_784 & _T_162; 
  assign _T_788 = _T_779 + _T_783; 
  assign _T_790 = _T_788 - _T_786; 
  assign _T_791 = _T_786 == 1'h0; 
  assign _T_793 = _T_791 | _T_779; 
  assign _T_795 = _T_793 | reset; 
  assign _T_796 = _T_795 == 1'h0; 
  assign _T_797 = _T_783 == 1'h0; 
  assign _T_798 = _T_779 != 1'h1; 
  assign _T_799 = _T_797 | _T_798; 
  assign _T_801 = _T_799 | reset; 
  assign _T_802 = _T_801 == 1'h0; 
  assign auto_in_a_ready = _T_68 & _T_71; 
  assign auto_in_d_valid = _T_87 ? auto_out_rvalid : auto_out_bvalid; 
  assign auto_in_d_bits_opcode = _T_87 ? 3'h1 : 3'h0; 
  assign auto_in_d_bits_size = _T_87 ? _T_46 : _T_48; 
  assign auto_in_d_bits_source = _T_87 ? _T_45 : _T_47; 
  assign auto_in_d_bits_denied = _T_87 ? _GEN_260 : _T_97; 
  assign auto_in_d_bits_data = auto_out_rdata; 
  assign auto_in_d_bits_corrupt = _T_87 ? _T_98 : 1'h0; 
  assign auto_out_awvalid = _T_52_valid & _T_52_bits_wen; 
  assign auto_out_awid = Queue_1_io_deq_bits_id; 
  assign auto_out_awaddr = Queue_1_io_deq_bits_addr; 
  assign auto_out_awlen = Queue_1_io_deq_bits_len; 
  assign auto_out_awsize = Queue_1_io_deq_bits_size; 
  assign auto_out_awburst = Queue_1_io_deq_bits_burst; 
  assign auto_out_awlock = Queue_1_io_deq_bits_lock; 
  assign auto_out_awcache = Queue_1_io_deq_bits_cache; 
  assign auto_out_awprot = Queue_1_io_deq_bits_prot; 
  assign auto_out_awqos = Queue_1_io_deq_bits_qos; 
  assign auto_out_awuser = Queue_1_io_deq_bits_user; 
  assign auto_out_awinstret = Queue_1_io_deq_bits_instret; 
  assign auto_out_wvalid = Queue_io_deq_valid; 
  assign auto_out_wdata = Queue_io_deq_bits_data; 
  assign auto_out_wstrb = Queue_io_deq_bits_strb; 
  assign auto_out_wlast = Queue_io_deq_bits_last; 
  assign auto_out_bready = auto_in_d_ready & _T_88; 
  assign auto_out_arvalid = _T_52_valid & _T_53; 
  assign auto_out_arid = Queue_1_io_deq_bits_id; 
  assign auto_out_araddr = Queue_1_io_deq_bits_addr; 
  assign auto_out_arlen = Queue_1_io_deq_bits_len; 
  assign auto_out_arsize = Queue_1_io_deq_bits_size; 
  assign auto_out_arburst = Queue_1_io_deq_bits_burst; 
  assign auto_out_arlock = Queue_1_io_deq_bits_lock; 
  assign auto_out_arcache = Queue_1_io_deq_bits_cache; 
  assign auto_out_arprot = Queue_1_io_deq_bits_prot; 
  assign auto_out_arqos = Queue_1_io_deq_bits_qos; 
  assign auto_out_aruser = Queue_1_io_deq_bits_user; 
  assign auto_out_arinstret = Queue_1_io_deq_bits_instret; 
  assign auto_out_rready = auto_in_d_ready; 
  assign TLMonitor_clock = clock; 
  assign TLMonitor_reset = reset; 
  assign TLMonitor_io_in_a_ready = _T_68 & _T_71; 
  assign TLMonitor_io_in_a_valid = auto_in_a_valid; 
  assign TLMonitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; 
  assign TLMonitor_io_in_a_bits_param = auto_in_a_bits_param; 
  assign TLMonitor_io_in_a_bits_size = auto_in_a_bits_size; 
  assign TLMonitor_io_in_a_bits_source = auto_in_a_bits_source; 
  assign TLMonitor_io_in_a_bits_address = auto_in_a_bits_address; 
  assign TLMonitor_io_in_a_bits_mask = auto_in_a_bits_mask; 
  assign TLMonitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; 
  assign TLMonitor_io_in_d_ready = auto_in_d_ready; 
  assign TLMonitor_io_in_d_valid = _T_87 ? auto_out_rvalid : auto_out_bvalid; 
  assign TLMonitor_io_in_d_bits_opcode = _T_87 ? 3'h1 : 3'h0; 
  assign TLMonitor_io_in_d_bits_size = _T_87 ? _T_46 : _T_48; 
  assign TLMonitor_io_in_d_bits_source = _T_87 ? _T_45 : _T_47; 
  assign TLMonitor_io_in_d_bits_denied = _T_87 ? _GEN_260 : _T_97; 
  assign TLMonitor_io_in_d_bits_corrupt = _T_87 ? _T_98 : 1'h0; 
  assign Queue_clock = clock; 
  assign Queue_reset = reset; 
  assign Queue_io_enq_valid = _T_81 & _T_69; 
  assign Queue_io_enq_bits_data = auto_in_a_bits_data; 
  assign Queue_io_enq_bits_strb = auto_in_a_bits_mask; 
  assign Queue_io_enq_bits_last = _T_27 | _T_28; 
  assign Queue_io_deq_ready = auto_out_wready; 
  assign Queue_1_clock = clock; 
  assign Queue_1_reset = reset; 
  assign Queue_1_io_enq_valid = _T_74 & _T_77; 
  assign Queue_1_io_enq_bits_id = 7'h7f == auto_in_a_bits_source ? 5'h6 : _GEN_128; 
  assign Queue_1_io_enq_bits_addr = auto_in_a_bits_address; 
  assign Queue_1_io_enq_bits_len = _T_63[10:3]; 
  assign Queue_1_io_enq_bits_size = _T_66[2:0]; 
  assign Queue_1_io_enq_bits_user = _GEN_284 | _T_43; 
  assign Queue_1_io_enq_bits_wen = _T_12 == 1'h0; 
  assign Queue_1_io_deq_ready = _T_52_bits_wen ? auto_out_awready : auto_out_arready; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_330 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_331 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_301 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_302 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_272 = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_273 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_243 = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_244 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_214 = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_215 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_185 = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_186 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_156 = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_157 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_779 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_751 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_723 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_695 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_667 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_639 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_611 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_583 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_555 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_527 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_499 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_471 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_443 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_415 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_387 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_359 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_23 = _RAND_30[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_57 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_84 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_91 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_94 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_330 <= 5'h0;
    end else begin
      _T_330 <= _T_341;
    end
    if (_T_334) begin
      _T_331 <= _T_13;
    end
    if (reset) begin
      _T_301 <= 5'h0;
    end else begin
      _T_301 <= _T_312;
    end
    if (_T_305) begin
      _T_302 <= _T_13;
    end
    if (reset) begin
      _T_272 <= 5'h0;
    end else begin
      _T_272 <= _T_283;
    end
    if (_T_276) begin
      _T_273 <= _T_13;
    end
    if (reset) begin
      _T_243 <= 5'h0;
    end else begin
      _T_243 <= _T_254;
    end
    if (_T_247) begin
      _T_244 <= _T_13;
    end
    if (reset) begin
      _T_214 <= 5'h0;
    end else begin
      _T_214 <= _T_225;
    end
    if (_T_218) begin
      _T_215 <= _T_13;
    end
    if (reset) begin
      _T_185 <= 5'h0;
    end else begin
      _T_185 <= _T_196;
    end
    if (_T_189) begin
      _T_186 <= _T_13;
    end
    if (reset) begin
      _T_156 <= 5'h0;
    end else begin
      _T_156 <= _T_167;
    end
    if (_T_160) begin
      _T_157 <= _T_13;
    end
    if (reset) begin
      _T_779 <= 1'h0;
    end else begin
      _T_779 <= _T_790;
    end
    if (reset) begin
      _T_751 <= 1'h0;
    end else begin
      _T_751 <= _T_762;
    end
    if (reset) begin
      _T_723 <= 1'h0;
    end else begin
      _T_723 <= _T_734;
    end
    if (reset) begin
      _T_695 <= 1'h0;
    end else begin
      _T_695 <= _T_706;
    end
    if (reset) begin
      _T_667 <= 1'h0;
    end else begin
      _T_667 <= _T_678;
    end
    if (reset) begin
      _T_639 <= 1'h0;
    end else begin
      _T_639 <= _T_650;
    end
    if (reset) begin
      _T_611 <= 1'h0;
    end else begin
      _T_611 <= _T_622;
    end
    if (reset) begin
      _T_583 <= 1'h0;
    end else begin
      _T_583 <= _T_594;
    end
    if (reset) begin
      _T_555 <= 1'h0;
    end else begin
      _T_555 <= _T_566;
    end
    if (reset) begin
      _T_527 <= 1'h0;
    end else begin
      _T_527 <= _T_538;
    end
    if (reset) begin
      _T_499 <= 1'h0;
    end else begin
      _T_499 <= _T_510;
    end
    if (reset) begin
      _T_471 <= 1'h0;
    end else begin
      _T_471 <= _T_482;
    end
    if (reset) begin
      _T_443 <= 1'h0;
    end else begin
      _T_443 <= _T_454;
    end
    if (reset) begin
      _T_415 <= 1'h0;
    end else begin
      _T_415 <= _T_426;
    end
    if (reset) begin
      _T_387 <= 1'h0;
    end else begin
      _T_387 <= _T_398;
    end
    if (reset) begin
      _T_359 <= 1'h0;
    end else begin
      _T_359 <= _T_370;
    end
    if (reset) begin
      _T_23 <= 5'h0;
    end else begin
      if (_T_14) begin
        if (_T_26) begin
          if (_T_13) begin
            _T_23 <= _T_19;
          end else begin
            _T_23 <= 5'h0;
          end
        end else begin
          _T_23 <= _T_25;
        end
      end
    end
    if (reset) begin
      _T_57 <= 1'h0;
    end else begin
      if (_T_14) begin
        _T_57 <= _T_59;
      end
    end
    if (reset) begin
      _T_84 <= 1'h0;
    end else begin
      if (_T_85) begin
        _T_84 <= _T_86;
      end
    end
    if (reset) begin
      _T_91 <= 1'h1;
    end else begin
      if (_T_85) begin
        _T_91 <= auto_out_rlast;
      end
    end
    if (_T_91) begin
      _T_94 <= _T_93;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:125 assert (a_source  < UInt(BigInt(1) << sourceBits))\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:126 assert (a_size    < UInt(BigInt(1) << sizeBits))\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_173) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_173) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_179) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_179) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_202) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_202) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_208) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_208) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_231) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_231) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_237) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_237) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_260) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_260) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_266) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_266) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_289) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_289) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_295) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_295) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_318) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_318) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_324) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_324) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_347) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_347) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_353) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_353) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_376) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_376) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_382) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_382) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_404) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_404) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_410) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_410) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_432) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_432) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_438) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_438) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_460) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_460) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_466) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_466) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_488) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_488) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_494) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_494) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_516) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_516) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_522) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_522) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_544) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_544) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_550) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_550) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_572) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_572) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_578) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_578) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_600) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_600) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_606) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_606) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_628) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_628) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_634) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_634) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_656) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_656) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_662) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_662) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_684) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_684) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_690) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_690) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_712) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_712) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_718) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_718) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_740) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_740) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_746) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_746) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_768) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_768) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_774) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_774) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_796) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_796) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_802) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_802) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLToAXI4( 
  input         clock, 
  input         reset, 
  output        auto_in_a_ready, 
  input         auto_in_a_valid, 
  input  [2:0]  auto_in_a_bits_opcode, 
  input  [2:0]  auto_in_a_bits_param, 
  input  [2:0]  auto_in_a_bits_size, 
  input  [6:0]  auto_in_a_bits_source, 
  input  [31:0] auto_in_a_bits_address, 
  input  [7:0]  auto_in_a_bits_mask, 
  input  [63:0] auto_in_a_bits_data, 
  input         auto_in_a_bits_corrupt, 
  input         auto_in_d_ready, 
  output        auto_in_d_valid, 
  output [2:0]  auto_in_d_bits_opcode, 
  output [2:0]  auto_in_d_bits_size, 
  output [6:0]  auto_in_d_bits_source, 
  output        auto_in_d_bits_denied, 
  output [63:0] auto_in_d_bits_data, 
  output        auto_in_d_bits_corrupt, 
  input         auto_out_awready, 
  output        auto_out_awvalid, 
  output [4:0]  auto_out_awid, 
  output [31:0] auto_out_awaddr, 
  output [7:0]  auto_out_awlen, 
  output [2:0]  auto_out_awsize, 
  output [1:0]  auto_out_awburst, 
  output        auto_out_awlock, 
  output [3:0]  auto_out_awcache, 
  output [2:0]  auto_out_awprot, 
  output [3:0]  auto_out_awqos, 
  output [10:0] auto_out_awuser, 
  output [63:0] auto_out_awinstret, 
  input         auto_out_wready, 
  output        auto_out_wvalid, 
  output [63:0] auto_out_wdata, 
  output [7:0]  auto_out_wstrb, 
  output        auto_out_wlast, 
  output        auto_out_bready, 
  input         auto_out_bvalid, 
  input  [4:0]  auto_out_bid, 
  input  [1:0]  auto_out_bresp, 
  input  [10:0] auto_out_buser, 
  input         auto_out_arready, 
  output        auto_out_arvalid, 
  output [4:0]  auto_out_arid, 
  output [31:0] auto_out_araddr, 
  output [7:0]  auto_out_arlen, 
  output [2:0]  auto_out_arsize, 
  output [1:0]  auto_out_arburst, 
  output        auto_out_arlock, 
  output [3:0]  auto_out_arcache, 
  output [2:0]  auto_out_arprot, 
  output [3:0]  auto_out_arqos, 
  output [10:0] auto_out_aruser, 
  output [63:0] auto_out_arinstret, 
  output        auto_out_rready, 
  input         auto_out_rvalid, 
  input  [4:0]  auto_out_rid, 
  input  [63:0] auto_out_rdata, 
  input  [1:0]  auto_out_rresp, 
  input  [10:0] auto_out_ruser, 
  input         auto_out_rlast 
);
  wire  TLMonitor_clock; 
  wire  TLMonitor_reset; 
  wire  TLMonitor_io_in_a_ready; 
  wire  TLMonitor_io_in_a_valid; 
  wire [2:0] TLMonitor_io_in_a_bits_opcode; 
  wire [2:0] TLMonitor_io_in_a_bits_param; 
  wire [2:0] TLMonitor_io_in_a_bits_size; 
  wire [6:0] TLMonitor_io_in_a_bits_source; 
  wire [31:0] TLMonitor_io_in_a_bits_address; 
  wire [7:0] TLMonitor_io_in_a_bits_mask; 
  wire  TLMonitor_io_in_a_bits_corrupt; 
  wire  TLMonitor_io_in_d_ready; 
  wire  TLMonitor_io_in_d_valid; 
  wire [2:0] TLMonitor_io_in_d_bits_opcode; 
  wire [2:0] TLMonitor_io_in_d_bits_size; 
  wire [6:0] TLMonitor_io_in_d_bits_source; 
  wire  TLMonitor_io_in_d_bits_denied; 
  wire  TLMonitor_io_in_d_bits_corrupt; 
  wire  Queue_clock; 
  wire  Queue_reset; 
  wire  Queue_io_enq_ready; 
  wire  Queue_io_enq_valid; 
  wire [63:0] Queue_io_enq_bits_data; 
  wire [7:0] Queue_io_enq_bits_strb; 
  wire  Queue_io_enq_bits_last; 
  wire  Queue_io_deq_ready; 
  wire  Queue_io_deq_valid; 
  wire [63:0] Queue_io_deq_bits_data; 
  wire [7:0] Queue_io_deq_bits_strb; 
  wire  Queue_io_deq_bits_last; 
  wire  Queue_1_clock; 
  wire  Queue_1_reset; 
  wire  Queue_1_io_enq_ready; 
  wire  Queue_1_io_enq_valid; 
  wire [4:0] Queue_1_io_enq_bits_id; 
  wire [31:0] Queue_1_io_enq_bits_addr; 
  wire [7:0] Queue_1_io_enq_bits_len; 
  wire [2:0] Queue_1_io_enq_bits_size; 
  wire [10:0] Queue_1_io_enq_bits_user; 
  wire  Queue_1_io_enq_bits_wen; 
  wire  Queue_1_io_deq_ready; 
  wire  Queue_1_io_deq_valid; 
  wire [4:0] Queue_1_io_deq_bits_id; 
  wire [31:0] Queue_1_io_deq_bits_addr; 
  wire [7:0] Queue_1_io_deq_bits_len; 
  wire [2:0] Queue_1_io_deq_bits_size; 
  wire [1:0] Queue_1_io_deq_bits_burst; 
  wire  Queue_1_io_deq_bits_lock; 
  wire [3:0] Queue_1_io_deq_bits_cache; 
  wire [2:0] Queue_1_io_deq_bits_prot; 
  wire [3:0] Queue_1_io_deq_bits_qos; 
  wire [10:0] Queue_1_io_deq_bits_user; 
  wire [63:0] Queue_1_io_deq_bits_instret; 
  wire  Queue_1_io_deq_bits_wen; 
  wire  _T_12; 
  wire  _T_13; 
  reg [4:0] _T_330; 
  reg [31:0] _RAND_0;
  wire  _T_332; 
  wire  _T_355; 
  reg  _T_331; 
  reg [31:0] _RAND_1;
  wire  _T_354; 
  wire  _T_356; 
  wire  _T_357; 
  wire  _T_358; 
  reg [4:0] _T_301; 
  reg [31:0] _RAND_2;
  wire  _T_303; 
  wire  _T_326; 
  reg  _T_302; 
  reg [31:0] _RAND_3;
  wire  _T_325; 
  wire  _T_327; 
  wire  _T_328; 
  wire  _T_329; 
  reg [4:0] _T_272; 
  reg [31:0] _RAND_4;
  wire  _T_274; 
  wire  _T_297; 
  reg  _T_273; 
  reg [31:0] _RAND_5;
  wire  _T_296; 
  wire  _T_298; 
  wire  _T_299; 
  wire  _T_300; 
  reg [4:0] _T_243; 
  reg [31:0] _RAND_6;
  wire  _T_245; 
  wire  _T_268; 
  reg  _T_244; 
  reg [31:0] _RAND_7;
  wire  _T_267; 
  wire  _T_269; 
  wire  _T_270; 
  wire  _T_271; 
  reg [4:0] _T_214; 
  reg [31:0] _RAND_8;
  wire  _T_216; 
  wire  _T_239; 
  reg  _T_215; 
  reg [31:0] _RAND_9;
  wire  _T_238; 
  wire  _T_240; 
  wire  _T_241; 
  wire  _T_242; 
  reg [4:0] _T_185; 
  reg [31:0] _RAND_10;
  wire  _T_187; 
  wire  _T_210; 
  reg  _T_186; 
  reg [31:0] _RAND_11;
  wire  _T_209; 
  wire  _T_211; 
  wire  _T_212; 
  wire  _T_213; 
  reg [4:0] _T_156; 
  reg [31:0] _RAND_12;
  wire  _T_158; 
  wire  _T_181; 
  reg  _T_157; 
  reg [31:0] _RAND_13;
  wire  _T_180; 
  wire  _T_182; 
  wire  _T_183; 
  wire  _T_184; 
  reg  _T_779; 
  reg [31:0] _RAND_14;
  reg  _T_751; 
  reg [31:0] _RAND_15;
  reg  _T_723; 
  reg [31:0] _RAND_16;
  reg  _T_695; 
  reg [31:0] _RAND_17;
  reg  _T_667; 
  reg [31:0] _RAND_18;
  reg  _T_639; 
  reg [31:0] _RAND_19;
  reg  _T_611; 
  reg [31:0] _RAND_20;
  reg  _T_583; 
  reg [31:0] _RAND_21;
  reg  _T_555; 
  reg [31:0] _RAND_22;
  reg  _T_527; 
  reg [31:0] _RAND_23;
  reg  _T_499; 
  reg [31:0] _RAND_24;
  reg  _T_471; 
  reg [31:0] _RAND_25;
  reg  _T_443; 
  reg [31:0] _RAND_26;
  reg  _T_415; 
  reg [31:0] _RAND_27;
  reg  _T_387; 
  reg [31:0] _RAND_28;
  reg  _T_359; 
  reg [31:0] _RAND_29;
  wire  _GEN_131; 
  wire  _GEN_132; 
  wire  _GEN_133; 
  wire  _GEN_134; 
  wire  _GEN_135; 
  wire  _GEN_136; 
  wire  _GEN_137; 
  wire  _GEN_138; 
  wire  _GEN_139; 
  wire  _GEN_140; 
  wire  _GEN_141; 
  wire  _GEN_142; 
  wire  _GEN_143; 
  wire  _GEN_144; 
  wire  _GEN_145; 
  wire  _GEN_146; 
  wire  _GEN_147; 
  wire  _GEN_148; 
  wire  _GEN_149; 
  wire  _GEN_150; 
  wire  _GEN_151; 
  wire  _GEN_152; 
  wire  _GEN_153; 
  wire  _GEN_154; 
  wire  _GEN_155; 
  wire  _GEN_156; 
  wire  _GEN_157; 
  wire  _GEN_158; 
  wire  _GEN_159; 
  wire  _GEN_160; 
  wire  _GEN_161; 
  wire  _GEN_162; 
  wire  _GEN_163; 
  wire  _GEN_164; 
  wire  _GEN_165; 
  wire  _GEN_166; 
  wire  _GEN_167; 
  wire  _GEN_168; 
  wire  _GEN_169; 
  wire  _GEN_170; 
  wire  _GEN_171; 
  wire  _GEN_172; 
  wire  _GEN_173; 
  wire  _GEN_174; 
  wire  _GEN_175; 
  wire  _GEN_176; 
  wire  _GEN_177; 
  wire  _GEN_178; 
  wire  _GEN_179; 
  wire  _GEN_180; 
  wire  _GEN_181; 
  wire  _GEN_182; 
  wire  _GEN_183; 
  wire  _GEN_184; 
  wire  _GEN_185; 
  wire  _GEN_186; 
  wire  _GEN_187; 
  wire  _GEN_188; 
  wire  _GEN_189; 
  wire  _GEN_190; 
  wire  _GEN_191; 
  wire  _GEN_192; 
  wire  _GEN_193; 
  wire  _GEN_194; 
  wire  _GEN_195; 
  wire  _GEN_196; 
  wire  _GEN_197; 
  wire  _GEN_198; 
  wire  _GEN_199; 
  wire  _GEN_200; 
  wire  _GEN_201; 
  wire  _GEN_202; 
  wire  _GEN_203; 
  wire  _GEN_204; 
  wire  _GEN_205; 
  wire  _GEN_206; 
  wire  _GEN_207; 
  wire  _GEN_208; 
  wire  _GEN_209; 
  wire  _GEN_210; 
  wire  _GEN_211; 
  wire  _GEN_212; 
  wire  _GEN_213; 
  wire  _GEN_214; 
  wire  _GEN_215; 
  wire  _GEN_216; 
  wire  _GEN_217; 
  wire  _GEN_218; 
  wire  _GEN_219; 
  wire  _GEN_220; 
  wire  _GEN_221; 
  wire  _GEN_222; 
  wire  _GEN_223; 
  wire  _GEN_224; 
  wire  _GEN_225; 
  wire  _GEN_226; 
  wire  _GEN_227; 
  wire  _GEN_228; 
  wire  _GEN_229; 
  wire  _GEN_230; 
  wire  _GEN_231; 
  wire  _GEN_232; 
  wire  _GEN_233; 
  wire  _GEN_234; 
  wire  _GEN_235; 
  wire  _GEN_236; 
  wire  _GEN_237; 
  wire  _GEN_238; 
  wire  _GEN_239; 
  wire  _GEN_240; 
  wire  _GEN_241; 
  wire  _GEN_242; 
  wire  _GEN_243; 
  wire  _GEN_244; 
  wire  _GEN_245; 
  wire  _GEN_246; 
  wire  _GEN_247; 
  wire  _GEN_248; 
  wire  _GEN_249; 
  wire  _GEN_250; 
  wire  _GEN_251; 
  wire  _GEN_252; 
  wire  _GEN_253; 
  wire  _GEN_254; 
  wire  _GEN_255; 
  wire  _GEN_256; 
  wire  _GEN_257; 
  reg [2:0] _T_23; 
  reg [31:0] _RAND_30;
  wire  _T_26; 
  wire  _T_67; 
  wire  _T_68; 
  reg  _T_57; 
  reg [31:0] _RAND_31;
  wire  _T_49_ready; 
  wire  _T_69; 
  wire  _T_50_ready; 
  wire  _T_70; 
  wire  _T_71; 
  wire  _T_72; 
  wire  _T_14; 
  wire [12:0] _T_16; 
  wire [5:0] _T_17; 
  wire [5:0] _T_18; 
  wire [2:0] _T_19; 
  wire [2:0] _T_22; 
  wire [2:0] _T_25; 
  wire  _T_27; 
  wire  _T_28; 
  wire  _T_29; 
  wire [9:0] _T_43; 
  wire [9:0] _GEN_284; 
  wire [9:0] _T_44; 
  wire [6:0] _T_45; 
  wire [2:0] _T_46; 
  wire [6:0] _T_47; 
  wire [2:0] _T_48; 
  wire  _T_52_bits_wen; 
  wire  _T_53; 
  wire  _T_52_valid; 
  wire  _T_59; 
  wire [4:0] _GEN_3; 
  wire [4:0] _GEN_4; 
  wire [4:0] _GEN_5; 
  wire [4:0] _GEN_6; 
  wire [4:0] _GEN_7; 
  wire [4:0] _GEN_8; 
  wire [4:0] _GEN_9; 
  wire [4:0] _GEN_10; 
  wire [4:0] _GEN_11; 
  wire [4:0] _GEN_12; 
  wire [4:0] _GEN_13; 
  wire [4:0] _GEN_14; 
  wire [4:0] _GEN_15; 
  wire [4:0] _GEN_16; 
  wire [4:0] _GEN_17; 
  wire [4:0] _GEN_18; 
  wire [4:0] _GEN_19; 
  wire [4:0] _GEN_20; 
  wire [4:0] _GEN_21; 
  wire [4:0] _GEN_22; 
  wire [4:0] _GEN_23; 
  wire [4:0] _GEN_24; 
  wire [4:0] _GEN_25; 
  wire [4:0] _GEN_26; 
  wire [4:0] _GEN_27; 
  wire [4:0] _GEN_28; 
  wire [4:0] _GEN_29; 
  wire [4:0] _GEN_30; 
  wire [4:0] _GEN_31; 
  wire [4:0] _GEN_32; 
  wire [4:0] _GEN_33; 
  wire [4:0] _GEN_34; 
  wire [4:0] _GEN_35; 
  wire [4:0] _GEN_36; 
  wire [4:0] _GEN_37; 
  wire [4:0] _GEN_38; 
  wire [4:0] _GEN_39; 
  wire [4:0] _GEN_40; 
  wire [4:0] _GEN_41; 
  wire [4:0] _GEN_42; 
  wire [4:0] _GEN_43; 
  wire [4:0] _GEN_44; 
  wire [4:0] _GEN_45; 
  wire [4:0] _GEN_46; 
  wire [4:0] _GEN_47; 
  wire [4:0] _GEN_48; 
  wire [4:0] _GEN_49; 
  wire [4:0] _GEN_50; 
  wire [4:0] _GEN_51; 
  wire [4:0] _GEN_52; 
  wire [4:0] _GEN_53; 
  wire [4:0] _GEN_54; 
  wire [4:0] _GEN_55; 
  wire [4:0] _GEN_56; 
  wire [4:0] _GEN_57; 
  wire [4:0] _GEN_58; 
  wire [4:0] _GEN_59; 
  wire [4:0] _GEN_60; 
  wire [4:0] _GEN_61; 
  wire [4:0] _GEN_62; 
  wire [4:0] _GEN_63; 
  wire [4:0] _GEN_64; 
  wire [4:0] _GEN_65; 
  wire [4:0] _GEN_66; 
  wire [4:0] _GEN_67; 
  wire [4:0] _GEN_68; 
  wire [4:0] _GEN_69; 
  wire [4:0] _GEN_70; 
  wire [4:0] _GEN_71; 
  wire [4:0] _GEN_72; 
  wire [4:0] _GEN_73; 
  wire [4:0] _GEN_74; 
  wire [4:0] _GEN_75; 
  wire [4:0] _GEN_76; 
  wire [4:0] _GEN_77; 
  wire [4:0] _GEN_78; 
  wire [4:0] _GEN_79; 
  wire [4:0] _GEN_80; 
  wire [4:0] _GEN_81; 
  wire [4:0] _GEN_82; 
  wire [4:0] _GEN_83; 
  wire [4:0] _GEN_84; 
  wire [4:0] _GEN_85; 
  wire [4:0] _GEN_86; 
  wire [4:0] _GEN_87; 
  wire [4:0] _GEN_88; 
  wire [4:0] _GEN_89; 
  wire [4:0] _GEN_90; 
  wire [4:0] _GEN_91; 
  wire [4:0] _GEN_92; 
  wire [4:0] _GEN_93; 
  wire [4:0] _GEN_94; 
  wire [4:0] _GEN_95; 
  wire [4:0] _GEN_96; 
  wire [4:0] _GEN_97; 
  wire [4:0] _GEN_98; 
  wire [4:0] _GEN_99; 
  wire [4:0] _GEN_100; 
  wire [4:0] _GEN_101; 
  wire [4:0] _GEN_102; 
  wire [4:0] _GEN_103; 
  wire [4:0] _GEN_104; 
  wire [4:0] _GEN_105; 
  wire [4:0] _GEN_106; 
  wire [4:0] _GEN_107; 
  wire [4:0] _GEN_108; 
  wire [4:0] _GEN_109; 
  wire [4:0] _GEN_110; 
  wire [4:0] _GEN_111; 
  wire [4:0] _GEN_112; 
  wire [4:0] _GEN_113; 
  wire [4:0] _GEN_114; 
  wire [4:0] _GEN_115; 
  wire [4:0] _GEN_116; 
  wire [4:0] _GEN_117; 
  wire [4:0] _GEN_118; 
  wire [4:0] _GEN_119; 
  wire [4:0] _GEN_120; 
  wire [4:0] _GEN_121; 
  wire [4:0] _GEN_122; 
  wire [4:0] _GEN_123; 
  wire [4:0] _GEN_124; 
  wire [4:0] _GEN_125; 
  wire [4:0] _GEN_126; 
  wire [4:0] _GEN_127; 
  wire [4:0] _GEN_128; 
  wire [4:0] _GEN_129; 
  wire [17:0] _T_61; 
  wire [10:0] _T_62; 
  wire [10:0] _T_63; 
  wire  _T_65; 
  wire  _T_74; 
  wire  _T_75; 
  wire  _T_76; 
  wire  _T_77; 
  wire  _T_78; 
  wire  _T_81; 
  reg  _T_84; 
  reg [31:0] _RAND_32;
  wire  _T_85; 
  wire  _T_86; 
  wire  _T_87; 
  wire  _T_88; 
  wire  _T_90; 
  reg  _T_91; 
  reg [31:0] _RAND_33;
  wire  _T_93; 
  reg  _T_94; 
  reg [31:0] _RAND_34;
  wire  _GEN_260; 
  wire  _T_96; 
  wire  _T_97; 
  wire  _T_98; 
  wire [31:0] _T_103; 
  wire [22:0] _T_104; 
  wire  _T_105; 
  wire  _T_106; 
  wire  _T_107; 
  wire  _T_108; 
  wire  _T_109; 
  wire  _T_110; 
  wire  _T_111; 
  wire  _T_112; 
  wire  _T_113; 
  wire  _T_114; 
  wire  _T_115; 
  wire  _T_116; 
  wire  _T_117; 
  wire  _T_118; 
  wire  _T_119; 
  wire  _T_120; 
  wire  _T_121; 
  wire  _T_122; 
  wire  _T_123; 
  wire  _T_124; 
  wire  _T_125; 
  wire  _T_126; 
  wire  _T_127; 
  wire [4:0] _T_128; 
  wire [31:0] _T_130; 
  wire [22:0] _T_131; 
  wire  _T_132; 
  wire  _T_133; 
  wire  _T_134; 
  wire  _T_135; 
  wire  _T_136; 
  wire  _T_137; 
  wire  _T_138; 
  wire  _T_139; 
  wire  _T_140; 
  wire  _T_141; 
  wire  _T_142; 
  wire  _T_143; 
  wire  _T_144; 
  wire  _T_145; 
  wire  _T_146; 
  wire  _T_147; 
  wire  _T_148; 
  wire  _T_149; 
  wire  _T_150; 
  wire  _T_151; 
  wire  _T_152; 
  wire  _T_153; 
  wire  _T_154; 
  wire  _T_155; 
  wire  _T_159; 
  wire  _T_160; 
  wire  _T_161; 
  wire  _T_162; 
  wire  _T_163; 
  wire [4:0] _GEN_285; 
  wire [4:0] _T_165; 
  wire [4:0] _GEN_286; 
  wire [4:0] _T_167; 
  wire  _T_168; 
  wire  _T_169; 
  wire  _T_170; 
  wire  _T_172; 
  wire  _T_173; 
  wire  _T_174; 
  wire  _T_175; 
  wire  _T_176; 
  wire  _T_178; 
  wire  _T_179; 
  wire  _T_189; 
  wire  _T_190; 
  wire  _T_192; 
  wire [4:0] _GEN_287; 
  wire [4:0] _T_194; 
  wire [4:0] _GEN_288; 
  wire [4:0] _T_196; 
  wire  _T_197; 
  wire  _T_198; 
  wire  _T_199; 
  wire  _T_201; 
  wire  _T_202; 
  wire  _T_203; 
  wire  _T_204; 
  wire  _T_205; 
  wire  _T_207; 
  wire  _T_208; 
  wire  _T_218; 
  wire  _T_219; 
  wire  _T_221; 
  wire [4:0] _GEN_289; 
  wire [4:0] _T_223; 
  wire [4:0] _GEN_290; 
  wire [4:0] _T_225; 
  wire  _T_226; 
  wire  _T_227; 
  wire  _T_228; 
  wire  _T_230; 
  wire  _T_231; 
  wire  _T_232; 
  wire  _T_233; 
  wire  _T_234; 
  wire  _T_236; 
  wire  _T_237; 
  wire  _T_247; 
  wire  _T_248; 
  wire  _T_250; 
  wire [4:0] _GEN_291; 
  wire [4:0] _T_252; 
  wire [4:0] _GEN_292; 
  wire [4:0] _T_254; 
  wire  _T_255; 
  wire  _T_256; 
  wire  _T_257; 
  wire  _T_259; 
  wire  _T_260; 
  wire  _T_261; 
  wire  _T_262; 
  wire  _T_263; 
  wire  _T_265; 
  wire  _T_266; 
  wire  _T_276; 
  wire  _T_277; 
  wire  _T_279; 
  wire [4:0] _GEN_293; 
  wire [4:0] _T_281; 
  wire [4:0] _GEN_294; 
  wire [4:0] _T_283; 
  wire  _T_284; 
  wire  _T_285; 
  wire  _T_286; 
  wire  _T_288; 
  wire  _T_289; 
  wire  _T_290; 
  wire  _T_291; 
  wire  _T_292; 
  wire  _T_294; 
  wire  _T_295; 
  wire  _T_305; 
  wire  _T_306; 
  wire  _T_308; 
  wire [4:0] _GEN_295; 
  wire [4:0] _T_310; 
  wire [4:0] _GEN_296; 
  wire [4:0] _T_312; 
  wire  _T_313; 
  wire  _T_314; 
  wire  _T_315; 
  wire  _T_317; 
  wire  _T_318; 
  wire  _T_319; 
  wire  _T_320; 
  wire  _T_321; 
  wire  _T_323; 
  wire  _T_324; 
  wire  _T_334; 
  wire  _T_335; 
  wire  _T_337; 
  wire [4:0] _GEN_297; 
  wire [4:0] _T_339; 
  wire [4:0] _GEN_298; 
  wire [4:0] _T_341; 
  wire  _T_342; 
  wire  _T_343; 
  wire  _T_344; 
  wire  _T_346; 
  wire  _T_347; 
  wire  _T_348; 
  wire  _T_349; 
  wire  _T_350; 
  wire  _T_352; 
  wire  _T_353; 
  wire  _T_363; 
  wire  _T_364; 
  wire  _T_366; 
  wire  _T_368; 
  wire  _T_370; 
  wire  _T_371; 
  wire  _T_373; 
  wire  _T_375; 
  wire  _T_376; 
  wire  _T_377; 
  wire  _T_378; 
  wire  _T_379; 
  wire  _T_381; 
  wire  _T_382; 
  wire  _T_391; 
  wire  _T_392; 
  wire  _T_394; 
  wire  _T_396; 
  wire  _T_398; 
  wire  _T_399; 
  wire  _T_401; 
  wire  _T_403; 
  wire  _T_404; 
  wire  _T_405; 
  wire  _T_406; 
  wire  _T_407; 
  wire  _T_409; 
  wire  _T_410; 
  wire  _T_419; 
  wire  _T_420; 
  wire  _T_422; 
  wire  _T_424; 
  wire  _T_426; 
  wire  _T_427; 
  wire  _T_429; 
  wire  _T_431; 
  wire  _T_432; 
  wire  _T_433; 
  wire  _T_434; 
  wire  _T_435; 
  wire  _T_437; 
  wire  _T_438; 
  wire  _T_447; 
  wire  _T_448; 
  wire  _T_450; 
  wire  _T_452; 
  wire  _T_454; 
  wire  _T_455; 
  wire  _T_457; 
  wire  _T_459; 
  wire  _T_460; 
  wire  _T_461; 
  wire  _T_462; 
  wire  _T_463; 
  wire  _T_465; 
  wire  _T_466; 
  wire  _T_475; 
  wire  _T_476; 
  wire  _T_478; 
  wire  _T_480; 
  wire  _T_482; 
  wire  _T_483; 
  wire  _T_485; 
  wire  _T_487; 
  wire  _T_488; 
  wire  _T_489; 
  wire  _T_490; 
  wire  _T_491; 
  wire  _T_493; 
  wire  _T_494; 
  wire  _T_503; 
  wire  _T_504; 
  wire  _T_506; 
  wire  _T_508; 
  wire  _T_510; 
  wire  _T_511; 
  wire  _T_513; 
  wire  _T_515; 
  wire  _T_516; 
  wire  _T_517; 
  wire  _T_518; 
  wire  _T_519; 
  wire  _T_521; 
  wire  _T_522; 
  wire  _T_531; 
  wire  _T_532; 
  wire  _T_534; 
  wire  _T_536; 
  wire  _T_538; 
  wire  _T_539; 
  wire  _T_541; 
  wire  _T_543; 
  wire  _T_544; 
  wire  _T_545; 
  wire  _T_546; 
  wire  _T_547; 
  wire  _T_549; 
  wire  _T_550; 
  wire  _T_559; 
  wire  _T_560; 
  wire  _T_562; 
  wire  _T_564; 
  wire  _T_566; 
  wire  _T_567; 
  wire  _T_569; 
  wire  _T_571; 
  wire  _T_572; 
  wire  _T_573; 
  wire  _T_574; 
  wire  _T_575; 
  wire  _T_577; 
  wire  _T_578; 
  wire  _T_587; 
  wire  _T_588; 
  wire  _T_590; 
  wire  _T_592; 
  wire  _T_594; 
  wire  _T_595; 
  wire  _T_597; 
  wire  _T_599; 
  wire  _T_600; 
  wire  _T_601; 
  wire  _T_602; 
  wire  _T_603; 
  wire  _T_605; 
  wire  _T_606; 
  wire  _T_615; 
  wire  _T_616; 
  wire  _T_618; 
  wire  _T_620; 
  wire  _T_622; 
  wire  _T_623; 
  wire  _T_625; 
  wire  _T_627; 
  wire  _T_628; 
  wire  _T_629; 
  wire  _T_630; 
  wire  _T_631; 
  wire  _T_633; 
  wire  _T_634; 
  wire  _T_643; 
  wire  _T_644; 
  wire  _T_646; 
  wire  _T_648; 
  wire  _T_650; 
  wire  _T_651; 
  wire  _T_653; 
  wire  _T_655; 
  wire  _T_656; 
  wire  _T_657; 
  wire  _T_658; 
  wire  _T_659; 
  wire  _T_661; 
  wire  _T_662; 
  wire  _T_671; 
  wire  _T_672; 
  wire  _T_674; 
  wire  _T_676; 
  wire  _T_678; 
  wire  _T_679; 
  wire  _T_681; 
  wire  _T_683; 
  wire  _T_684; 
  wire  _T_685; 
  wire  _T_686; 
  wire  _T_687; 
  wire  _T_689; 
  wire  _T_690; 
  wire  _T_699; 
  wire  _T_700; 
  wire  _T_702; 
  wire  _T_704; 
  wire  _T_706; 
  wire  _T_707; 
  wire  _T_709; 
  wire  _T_711; 
  wire  _T_712; 
  wire  _T_713; 
  wire  _T_714; 
  wire  _T_715; 
  wire  _T_717; 
  wire  _T_718; 
  wire  _T_727; 
  wire  _T_728; 
  wire  _T_730; 
  wire  _T_732; 
  wire  _T_734; 
  wire  _T_735; 
  wire  _T_737; 
  wire  _T_739; 
  wire  _T_740; 
  wire  _T_741; 
  wire  _T_742; 
  wire  _T_743; 
  wire  _T_745; 
  wire  _T_746; 
  wire  _T_755; 
  wire  _T_756; 
  wire  _T_758; 
  wire  _T_760; 
  wire  _T_762; 
  wire  _T_763; 
  wire  _T_765; 
  wire  _T_767; 
  wire  _T_768; 
  wire  _T_769; 
  wire  _T_770; 
  wire  _T_771; 
  wire  _T_773; 
  wire  _T_774; 
  wire  _T_783; 
  wire  _T_784; 
  wire  _T_786; 
  wire  _T_788; 
  wire  _T_790; 
  wire  _T_791; 
  wire  _T_793; 
  wire  _T_795; 
  wire  _T_796; 
  wire  _T_797; 
  wire  _T_798; 
  wire  _T_799; 
  wire  _T_801; 
  wire  _T_802; 
  dual_TLMonitor_9 dual_TLMonitor ( 
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_io_in_a_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt)
  );
  dual_Queue_46 dual_Queue ( 
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_strb(Queue_io_enq_bits_strb),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_strb(Queue_io_deq_bits_strb),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  dual_Queue_47 Queue_1 ( 
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_id(Queue_1_io_enq_bits_id),
    .io_enq_bits_addr(Queue_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_user(Queue_1_io_enq_bits_user),
    .io_enq_bits_wen(Queue_1_io_enq_bits_wen),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_id(Queue_1_io_deq_bits_id),
    .io_deq_bits_addr(Queue_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_1_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_1_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_1_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_1_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_1_io_deq_bits_qos),
    .io_deq_bits_user(Queue_1_io_deq_bits_user),
    .io_deq_bits_instret(Queue_1_io_deq_bits_instret),
    .io_deq_bits_wen(Queue_1_io_deq_bits_wen)
  );
  assign _T_12 = auto_in_a_bits_opcode[2]; 
  assign _T_13 = _T_12 == 1'h0; 
  assign _T_332 = _T_330 == 5'h0; 
  assign _T_355 = _T_332 == 1'h0; 
  assign _T_354 = _T_331 != _T_13; 
  assign _T_356 = _T_355 & _T_354; 
  assign _T_357 = _T_330 == 5'h10; 
  assign _T_358 = _T_356 | _T_357; 
  assign _T_303 = _T_301 == 5'h0; 
  assign _T_326 = _T_303 == 1'h0; 
  assign _T_325 = _T_302 != _T_13; 
  assign _T_327 = _T_326 & _T_325; 
  assign _T_328 = _T_301 == 5'h10; 
  assign _T_329 = _T_327 | _T_328; 
  assign _T_274 = _T_272 == 5'h0; 
  assign _T_297 = _T_274 == 1'h0; 
  assign _T_296 = _T_273 != _T_13; 
  assign _T_298 = _T_297 & _T_296; 
  assign _T_299 = _T_272 == 5'h10; 
  assign _T_300 = _T_298 | _T_299; 
  assign _T_245 = _T_243 == 5'h0; 
  assign _T_268 = _T_245 == 1'h0; 
  assign _T_267 = _T_244 != _T_13; 
  assign _T_269 = _T_268 & _T_267; 
  assign _T_270 = _T_243 == 5'h10; 
  assign _T_271 = _T_269 | _T_270; 
  assign _T_216 = _T_214 == 5'h0; 
  assign _T_239 = _T_216 == 1'h0; 
  assign _T_238 = _T_215 != _T_13; 
  assign _T_240 = _T_239 & _T_238; 
  assign _T_241 = _T_214 == 5'h10; 
  assign _T_242 = _T_240 | _T_241; 
  assign _T_187 = _T_185 == 5'h0; 
  assign _T_210 = _T_187 == 1'h0; 
  assign _T_209 = _T_186 != _T_13; 
  assign _T_211 = _T_210 & _T_209; 
  assign _T_212 = _T_185 == 5'h10; 
  assign _T_213 = _T_211 | _T_212; 
  assign _T_158 = _T_156 == 5'h0; 
  assign _T_181 = _T_158 == 1'h0; 
  assign _T_180 = _T_157 != _T_13; 
  assign _T_182 = _T_181 & _T_180; 
  assign _T_183 = _T_156 == 5'h10; 
  assign _T_184 = _T_182 | _T_183; 
  assign _GEN_131 = 7'h1 == auto_in_a_bits_source ? _T_387 : _T_359; 
  assign _GEN_132 = 7'h2 == auto_in_a_bits_source ? _T_415 : _GEN_131; 
  assign _GEN_133 = 7'h3 == auto_in_a_bits_source ? _T_443 : _GEN_132; 
  assign _GEN_134 = 7'h4 == auto_in_a_bits_source ? _T_471 : _GEN_133; 
  assign _GEN_135 = 7'h5 == auto_in_a_bits_source ? _T_499 : _GEN_134; 
  assign _GEN_136 = 7'h6 == auto_in_a_bits_source ? _T_527 : _GEN_135; 
  assign _GEN_137 = 7'h7 == auto_in_a_bits_source ? _T_555 : _GEN_136; 
  assign _GEN_138 = 7'h8 == auto_in_a_bits_source ? _T_583 : _GEN_137; 
  assign _GEN_139 = 7'h9 == auto_in_a_bits_source ? _T_611 : _GEN_138; 
  assign _GEN_140 = 7'ha == auto_in_a_bits_source ? _T_639 : _GEN_139; 
  assign _GEN_141 = 7'hb == auto_in_a_bits_source ? _T_667 : _GEN_140; 
  assign _GEN_142 = 7'hc == auto_in_a_bits_source ? _T_695 : _GEN_141; 
  assign _GEN_143 = 7'hd == auto_in_a_bits_source ? _T_723 : _GEN_142; 
  assign _GEN_144 = 7'he == auto_in_a_bits_source ? _T_751 : _GEN_143; 
  assign _GEN_145 = 7'hf == auto_in_a_bits_source ? _T_779 : _GEN_144; 
  assign _GEN_146 = 7'h10 == auto_in_a_bits_source ? _T_184 : _GEN_145; 
  assign _GEN_147 = 7'h11 == auto_in_a_bits_source ? _T_184 : _GEN_146; 
  assign _GEN_148 = 7'h12 == auto_in_a_bits_source ? _T_184 : _GEN_147; 
  assign _GEN_149 = 7'h13 == auto_in_a_bits_source ? _T_184 : _GEN_148; 
  assign _GEN_150 = 7'h14 == auto_in_a_bits_source ? _T_184 : _GEN_149; 
  assign _GEN_151 = 7'h15 == auto_in_a_bits_source ? _T_184 : _GEN_150; 
  assign _GEN_152 = 7'h16 == auto_in_a_bits_source ? _T_184 : _GEN_151; 
  assign _GEN_153 = 7'h17 == auto_in_a_bits_source ? _T_184 : _GEN_152; 
  assign _GEN_154 = 7'h18 == auto_in_a_bits_source ? _T_184 : _GEN_153; 
  assign _GEN_155 = 7'h19 == auto_in_a_bits_source ? _T_184 : _GEN_154; 
  assign _GEN_156 = 7'h1a == auto_in_a_bits_source ? _T_184 : _GEN_155; 
  assign _GEN_157 = 7'h1b == auto_in_a_bits_source ? _T_184 : _GEN_156; 
  assign _GEN_158 = 7'h1c == auto_in_a_bits_source ? _T_184 : _GEN_157; 
  assign _GEN_159 = 7'h1d == auto_in_a_bits_source ? _T_184 : _GEN_158; 
  assign _GEN_160 = 7'h1e == auto_in_a_bits_source ? _T_184 : _GEN_159; 
  assign _GEN_161 = 7'h1f == auto_in_a_bits_source ? _T_184 : _GEN_160; 
  assign _GEN_162 = 7'h20 == auto_in_a_bits_source ? _T_213 : _GEN_161; 
  assign _GEN_163 = 7'h21 == auto_in_a_bits_source ? _T_213 : _GEN_162; 
  assign _GEN_164 = 7'h22 == auto_in_a_bits_source ? _T_213 : _GEN_163; 
  assign _GEN_165 = 7'h23 == auto_in_a_bits_source ? _T_213 : _GEN_164; 
  assign _GEN_166 = 7'h24 == auto_in_a_bits_source ? _T_213 : _GEN_165; 
  assign _GEN_167 = 7'h25 == auto_in_a_bits_source ? _T_213 : _GEN_166; 
  assign _GEN_168 = 7'h26 == auto_in_a_bits_source ? _T_213 : _GEN_167; 
  assign _GEN_169 = 7'h27 == auto_in_a_bits_source ? _T_213 : _GEN_168; 
  assign _GEN_170 = 7'h28 == auto_in_a_bits_source ? _T_213 : _GEN_169; 
  assign _GEN_171 = 7'h29 == auto_in_a_bits_source ? _T_213 : _GEN_170; 
  assign _GEN_172 = 7'h2a == auto_in_a_bits_source ? _T_213 : _GEN_171; 
  assign _GEN_173 = 7'h2b == auto_in_a_bits_source ? _T_213 : _GEN_172; 
  assign _GEN_174 = 7'h2c == auto_in_a_bits_source ? _T_213 : _GEN_173; 
  assign _GEN_175 = 7'h2d == auto_in_a_bits_source ? _T_213 : _GEN_174; 
  assign _GEN_176 = 7'h2e == auto_in_a_bits_source ? _T_213 : _GEN_175; 
  assign _GEN_177 = 7'h2f == auto_in_a_bits_source ? _T_213 : _GEN_176; 
  assign _GEN_178 = 7'h30 == auto_in_a_bits_source ? _T_242 : _GEN_177; 
  assign _GEN_179 = 7'h31 == auto_in_a_bits_source ? _T_242 : _GEN_178; 
  assign _GEN_180 = 7'h32 == auto_in_a_bits_source ? _T_242 : _GEN_179; 
  assign _GEN_181 = 7'h33 == auto_in_a_bits_source ? _T_242 : _GEN_180; 
  assign _GEN_182 = 7'h34 == auto_in_a_bits_source ? _T_242 : _GEN_181; 
  assign _GEN_183 = 7'h35 == auto_in_a_bits_source ? _T_242 : _GEN_182; 
  assign _GEN_184 = 7'h36 == auto_in_a_bits_source ? _T_242 : _GEN_183; 
  assign _GEN_185 = 7'h37 == auto_in_a_bits_source ? _T_242 : _GEN_184; 
  assign _GEN_186 = 7'h38 == auto_in_a_bits_source ? _T_242 : _GEN_185; 
  assign _GEN_187 = 7'h39 == auto_in_a_bits_source ? _T_242 : _GEN_186; 
  assign _GEN_188 = 7'h3a == auto_in_a_bits_source ? _T_242 : _GEN_187; 
  assign _GEN_189 = 7'h3b == auto_in_a_bits_source ? _T_242 : _GEN_188; 
  assign _GEN_190 = 7'h3c == auto_in_a_bits_source ? _T_242 : _GEN_189; 
  assign _GEN_191 = 7'h3d == auto_in_a_bits_source ? _T_242 : _GEN_190; 
  assign _GEN_192 = 7'h3e == auto_in_a_bits_source ? _T_242 : _GEN_191; 
  assign _GEN_193 = 7'h3f == auto_in_a_bits_source ? _T_242 : _GEN_192; 
  assign _GEN_194 = 7'h40 == auto_in_a_bits_source ? _T_271 : _GEN_193; 
  assign _GEN_195 = 7'h41 == auto_in_a_bits_source ? _T_271 : _GEN_194; 
  assign _GEN_196 = 7'h42 == auto_in_a_bits_source ? _T_271 : _GEN_195; 
  assign _GEN_197 = 7'h43 == auto_in_a_bits_source ? _T_271 : _GEN_196; 
  assign _GEN_198 = 7'h44 == auto_in_a_bits_source ? _T_271 : _GEN_197; 
  assign _GEN_199 = 7'h45 == auto_in_a_bits_source ? _T_271 : _GEN_198; 
  assign _GEN_200 = 7'h46 == auto_in_a_bits_source ? _T_271 : _GEN_199; 
  assign _GEN_201 = 7'h47 == auto_in_a_bits_source ? _T_271 : _GEN_200; 
  assign _GEN_202 = 7'h48 == auto_in_a_bits_source ? _T_271 : _GEN_201; 
  assign _GEN_203 = 7'h49 == auto_in_a_bits_source ? _T_271 : _GEN_202; 
  assign _GEN_204 = 7'h4a == auto_in_a_bits_source ? _T_271 : _GEN_203; 
  assign _GEN_205 = 7'h4b == auto_in_a_bits_source ? _T_271 : _GEN_204; 
  assign _GEN_206 = 7'h4c == auto_in_a_bits_source ? _T_271 : _GEN_205; 
  assign _GEN_207 = 7'h4d == auto_in_a_bits_source ? _T_271 : _GEN_206; 
  assign _GEN_208 = 7'h4e == auto_in_a_bits_source ? _T_271 : _GEN_207; 
  assign _GEN_209 = 7'h4f == auto_in_a_bits_source ? _T_271 : _GEN_208; 
  assign _GEN_210 = 7'h50 == auto_in_a_bits_source ? _T_300 : _GEN_209; 
  assign _GEN_211 = 7'h51 == auto_in_a_bits_source ? _T_300 : _GEN_210; 
  assign _GEN_212 = 7'h52 == auto_in_a_bits_source ? _T_300 : _GEN_211; 
  assign _GEN_213 = 7'h53 == auto_in_a_bits_source ? _T_300 : _GEN_212; 
  assign _GEN_214 = 7'h54 == auto_in_a_bits_source ? _T_300 : _GEN_213; 
  assign _GEN_215 = 7'h55 == auto_in_a_bits_source ? _T_300 : _GEN_214; 
  assign _GEN_216 = 7'h56 == auto_in_a_bits_source ? _T_300 : _GEN_215; 
  assign _GEN_217 = 7'h57 == auto_in_a_bits_source ? _T_300 : _GEN_216; 
  assign _GEN_218 = 7'h58 == auto_in_a_bits_source ? _T_300 : _GEN_217; 
  assign _GEN_219 = 7'h59 == auto_in_a_bits_source ? _T_300 : _GEN_218; 
  assign _GEN_220 = 7'h5a == auto_in_a_bits_source ? _T_300 : _GEN_219; 
  assign _GEN_221 = 7'h5b == auto_in_a_bits_source ? _T_300 : _GEN_220; 
  assign _GEN_222 = 7'h5c == auto_in_a_bits_source ? _T_300 : _GEN_221; 
  assign _GEN_223 = 7'h5d == auto_in_a_bits_source ? _T_300 : _GEN_222; 
  assign _GEN_224 = 7'h5e == auto_in_a_bits_source ? _T_300 : _GEN_223; 
  assign _GEN_225 = 7'h5f == auto_in_a_bits_source ? _T_300 : _GEN_224; 
  assign _GEN_226 = 7'h60 == auto_in_a_bits_source ? _T_329 : _GEN_225; 
  assign _GEN_227 = 7'h61 == auto_in_a_bits_source ? _T_329 : _GEN_226; 
  assign _GEN_228 = 7'h62 == auto_in_a_bits_source ? _T_329 : _GEN_227; 
  assign _GEN_229 = 7'h63 == auto_in_a_bits_source ? _T_329 : _GEN_228; 
  assign _GEN_230 = 7'h64 == auto_in_a_bits_source ? _T_329 : _GEN_229; 
  assign _GEN_231 = 7'h65 == auto_in_a_bits_source ? _T_329 : _GEN_230; 
  assign _GEN_232 = 7'h66 == auto_in_a_bits_source ? _T_329 : _GEN_231; 
  assign _GEN_233 = 7'h67 == auto_in_a_bits_source ? _T_329 : _GEN_232; 
  assign _GEN_234 = 7'h68 == auto_in_a_bits_source ? _T_329 : _GEN_233; 
  assign _GEN_235 = 7'h69 == auto_in_a_bits_source ? _T_329 : _GEN_234; 
  assign _GEN_236 = 7'h6a == auto_in_a_bits_source ? _T_329 : _GEN_235; 
  assign _GEN_237 = 7'h6b == auto_in_a_bits_source ? _T_329 : _GEN_236; 
  assign _GEN_238 = 7'h6c == auto_in_a_bits_source ? _T_329 : _GEN_237; 
  assign _GEN_239 = 7'h6d == auto_in_a_bits_source ? _T_329 : _GEN_238; 
  assign _GEN_240 = 7'h6e == auto_in_a_bits_source ? _T_329 : _GEN_239; 
  assign _GEN_241 = 7'h6f == auto_in_a_bits_source ? _T_329 : _GEN_240; 
  assign _GEN_242 = 7'h70 == auto_in_a_bits_source ? _T_358 : _GEN_241; 
  assign _GEN_243 = 7'h71 == auto_in_a_bits_source ? _T_358 : _GEN_242; 
  assign _GEN_244 = 7'h72 == auto_in_a_bits_source ? _T_358 : _GEN_243; 
  assign _GEN_245 = 7'h73 == auto_in_a_bits_source ? _T_358 : _GEN_244; 
  assign _GEN_246 = 7'h74 == auto_in_a_bits_source ? _T_358 : _GEN_245; 
  assign _GEN_247 = 7'h75 == auto_in_a_bits_source ? _T_358 : _GEN_246; 
  assign _GEN_248 = 7'h76 == auto_in_a_bits_source ? _T_358 : _GEN_247; 
  assign _GEN_249 = 7'h77 == auto_in_a_bits_source ? _T_358 : _GEN_248; 
  assign _GEN_250 = 7'h78 == auto_in_a_bits_source ? _T_358 : _GEN_249; 
  assign _GEN_251 = 7'h79 == auto_in_a_bits_source ? _T_358 : _GEN_250; 
  assign _GEN_252 = 7'h7a == auto_in_a_bits_source ? _T_358 : _GEN_251; 
  assign _GEN_253 = 7'h7b == auto_in_a_bits_source ? _T_358 : _GEN_252; 
  assign _GEN_254 = 7'h7c == auto_in_a_bits_source ? _T_358 : _GEN_253; 
  assign _GEN_255 = 7'h7d == auto_in_a_bits_source ? _T_358 : _GEN_254; 
  assign _GEN_256 = 7'h7e == auto_in_a_bits_source ? _T_358 : _GEN_255; 
  assign _GEN_257 = 7'h7f == auto_in_a_bits_source ? _T_358 : _GEN_256; 
  assign _T_26 = _T_23 == 3'h0; 
  assign _T_67 = _GEN_257 & _T_26; 
  assign _T_68 = _T_67 == 1'h0; 
  assign _T_49_ready = Queue_1_io_enq_ready; 
  assign _T_69 = _T_57 | _T_49_ready; 
  assign _T_50_ready = Queue_io_enq_ready; 
  assign _T_70 = _T_69 & _T_50_ready; 
  assign _T_71 = _T_13 ? _T_70 : _T_49_ready; 
  assign _T_72 = _T_68 & _T_71; 
  assign _T_14 = _T_72 & auto_in_a_valid; 
  assign _T_16 = 13'h3f << auto_in_a_bits_size; 
  assign _T_17 = _T_16[5:0]; 
  assign _T_18 = ~ _T_17; 
  assign _T_19 = _T_18[5:3]; 
  assign _T_22 = _T_13 ? _T_19 : 3'h0; 
  assign _T_25 = _T_23 - 3'h1; 
  assign _T_27 = _T_23 == 3'h1; 
  assign _T_28 = _T_22 == 3'h0; 
  assign _T_29 = _T_27 | _T_28; 
  assign _T_43 = {auto_in_a_bits_size, 7'h0}; 
  assign _GEN_284 = {{3'd0}, auto_in_a_bits_source}; 
  assign _T_44 = _GEN_284 | _T_43; 
  assign _T_45 = auto_out_ruser[6:0]; 
  assign _T_46 = auto_out_ruser[9:7]; 
  assign _T_47 = auto_out_buser[6:0]; 
  assign _T_48 = auto_out_buser[9:7]; 
  assign _T_52_bits_wen = Queue_1_io_deq_bits_wen; 
  assign _T_53 = _T_52_bits_wen == 1'h0; 
  assign _T_52_valid = Queue_1_io_deq_valid; 
  assign _T_59 = _T_29 == 1'h0; 
  assign _GEN_3 = 7'h1 == auto_in_a_bits_source ? 5'h8 : 5'h7; 
  assign _GEN_4 = 7'h2 == auto_in_a_bits_source ? 5'h9 : _GEN_3; 
  assign _GEN_5 = 7'h3 == auto_in_a_bits_source ? 5'ha : _GEN_4; 
  assign _GEN_6 = 7'h4 == auto_in_a_bits_source ? 5'hb : _GEN_5; 
  assign _GEN_7 = 7'h5 == auto_in_a_bits_source ? 5'hc : _GEN_6; 
  assign _GEN_8 = 7'h6 == auto_in_a_bits_source ? 5'hd : _GEN_7; 
  assign _GEN_9 = 7'h7 == auto_in_a_bits_source ? 5'he : _GEN_8; 
  assign _GEN_10 = 7'h8 == auto_in_a_bits_source ? 5'hf : _GEN_9; 
  assign _GEN_11 = 7'h9 == auto_in_a_bits_source ? 5'h10 : _GEN_10; 
  assign _GEN_12 = 7'ha == auto_in_a_bits_source ? 5'h11 : _GEN_11; 
  assign _GEN_13 = 7'hb == auto_in_a_bits_source ? 5'h12 : _GEN_12; 
  assign _GEN_14 = 7'hc == auto_in_a_bits_source ? 5'h13 : _GEN_13; 
  assign _GEN_15 = 7'hd == auto_in_a_bits_source ? 5'h14 : _GEN_14; 
  assign _GEN_16 = 7'he == auto_in_a_bits_source ? 5'h15 : _GEN_15; 
  assign _GEN_17 = 7'hf == auto_in_a_bits_source ? 5'h16 : _GEN_16; 
  assign _GEN_18 = 7'h10 == auto_in_a_bits_source ? 5'h0 : _GEN_17; 
  assign _GEN_19 = 7'h11 == auto_in_a_bits_source ? 5'h0 : _GEN_18; 
  assign _GEN_20 = 7'h12 == auto_in_a_bits_source ? 5'h0 : _GEN_19; 
  assign _GEN_21 = 7'h13 == auto_in_a_bits_source ? 5'h0 : _GEN_20; 
  assign _GEN_22 = 7'h14 == auto_in_a_bits_source ? 5'h0 : _GEN_21; 
  assign _GEN_23 = 7'h15 == auto_in_a_bits_source ? 5'h0 : _GEN_22; 
  assign _GEN_24 = 7'h16 == auto_in_a_bits_source ? 5'h0 : _GEN_23; 
  assign _GEN_25 = 7'h17 == auto_in_a_bits_source ? 5'h0 : _GEN_24; 
  assign _GEN_26 = 7'h18 == auto_in_a_bits_source ? 5'h0 : _GEN_25; 
  assign _GEN_27 = 7'h19 == auto_in_a_bits_source ? 5'h0 : _GEN_26; 
  assign _GEN_28 = 7'h1a == auto_in_a_bits_source ? 5'h0 : _GEN_27; 
  assign _GEN_29 = 7'h1b == auto_in_a_bits_source ? 5'h0 : _GEN_28; 
  assign _GEN_30 = 7'h1c == auto_in_a_bits_source ? 5'h0 : _GEN_29; 
  assign _GEN_31 = 7'h1d == auto_in_a_bits_source ? 5'h0 : _GEN_30; 
  assign _GEN_32 = 7'h1e == auto_in_a_bits_source ? 5'h0 : _GEN_31; 
  assign _GEN_33 = 7'h1f == auto_in_a_bits_source ? 5'h0 : _GEN_32; 
  assign _GEN_34 = 7'h20 == auto_in_a_bits_source ? 5'h1 : _GEN_33; 
  assign _GEN_35 = 7'h21 == auto_in_a_bits_source ? 5'h1 : _GEN_34; 
  assign _GEN_36 = 7'h22 == auto_in_a_bits_source ? 5'h1 : _GEN_35; 
  assign _GEN_37 = 7'h23 == auto_in_a_bits_source ? 5'h1 : _GEN_36; 
  assign _GEN_38 = 7'h24 == auto_in_a_bits_source ? 5'h1 : _GEN_37; 
  assign _GEN_39 = 7'h25 == auto_in_a_bits_source ? 5'h1 : _GEN_38; 
  assign _GEN_40 = 7'h26 == auto_in_a_bits_source ? 5'h1 : _GEN_39; 
  assign _GEN_41 = 7'h27 == auto_in_a_bits_source ? 5'h1 : _GEN_40; 
  assign _GEN_42 = 7'h28 == auto_in_a_bits_source ? 5'h1 : _GEN_41; 
  assign _GEN_43 = 7'h29 == auto_in_a_bits_source ? 5'h1 : _GEN_42; 
  assign _GEN_44 = 7'h2a == auto_in_a_bits_source ? 5'h1 : _GEN_43; 
  assign _GEN_45 = 7'h2b == auto_in_a_bits_source ? 5'h1 : _GEN_44; 
  assign _GEN_46 = 7'h2c == auto_in_a_bits_source ? 5'h1 : _GEN_45; 
  assign _GEN_47 = 7'h2d == auto_in_a_bits_source ? 5'h1 : _GEN_46; 
  assign _GEN_48 = 7'h2e == auto_in_a_bits_source ? 5'h1 : _GEN_47; 
  assign _GEN_49 = 7'h2f == auto_in_a_bits_source ? 5'h1 : _GEN_48; 
  assign _GEN_50 = 7'h30 == auto_in_a_bits_source ? 5'h2 : _GEN_49; 
  assign _GEN_51 = 7'h31 == auto_in_a_bits_source ? 5'h2 : _GEN_50; 
  assign _GEN_52 = 7'h32 == auto_in_a_bits_source ? 5'h2 : _GEN_51; 
  assign _GEN_53 = 7'h33 == auto_in_a_bits_source ? 5'h2 : _GEN_52; 
  assign _GEN_54 = 7'h34 == auto_in_a_bits_source ? 5'h2 : _GEN_53; 
  assign _GEN_55 = 7'h35 == auto_in_a_bits_source ? 5'h2 : _GEN_54; 
  assign _GEN_56 = 7'h36 == auto_in_a_bits_source ? 5'h2 : _GEN_55; 
  assign _GEN_57 = 7'h37 == auto_in_a_bits_source ? 5'h2 : _GEN_56; 
  assign _GEN_58 = 7'h38 == auto_in_a_bits_source ? 5'h2 : _GEN_57; 
  assign _GEN_59 = 7'h39 == auto_in_a_bits_source ? 5'h2 : _GEN_58; 
  assign _GEN_60 = 7'h3a == auto_in_a_bits_source ? 5'h2 : _GEN_59; 
  assign _GEN_61 = 7'h3b == auto_in_a_bits_source ? 5'h2 : _GEN_60; 
  assign _GEN_62 = 7'h3c == auto_in_a_bits_source ? 5'h2 : _GEN_61; 
  assign _GEN_63 = 7'h3d == auto_in_a_bits_source ? 5'h2 : _GEN_62; 
  assign _GEN_64 = 7'h3e == auto_in_a_bits_source ? 5'h2 : _GEN_63; 
  assign _GEN_65 = 7'h3f == auto_in_a_bits_source ? 5'h2 : _GEN_64; 
  assign _GEN_66 = 7'h40 == auto_in_a_bits_source ? 5'h3 : _GEN_65; 
  assign _GEN_67 = 7'h41 == auto_in_a_bits_source ? 5'h3 : _GEN_66; 
  assign _GEN_68 = 7'h42 == auto_in_a_bits_source ? 5'h3 : _GEN_67; 
  assign _GEN_69 = 7'h43 == auto_in_a_bits_source ? 5'h3 : _GEN_68; 
  assign _GEN_70 = 7'h44 == auto_in_a_bits_source ? 5'h3 : _GEN_69; 
  assign _GEN_71 = 7'h45 == auto_in_a_bits_source ? 5'h3 : _GEN_70; 
  assign _GEN_72 = 7'h46 == auto_in_a_bits_source ? 5'h3 : _GEN_71; 
  assign _GEN_73 = 7'h47 == auto_in_a_bits_source ? 5'h3 : _GEN_72; 
  assign _GEN_74 = 7'h48 == auto_in_a_bits_source ? 5'h3 : _GEN_73; 
  assign _GEN_75 = 7'h49 == auto_in_a_bits_source ? 5'h3 : _GEN_74; 
  assign _GEN_76 = 7'h4a == auto_in_a_bits_source ? 5'h3 : _GEN_75; 
  assign _GEN_77 = 7'h4b == auto_in_a_bits_source ? 5'h3 : _GEN_76; 
  assign _GEN_78 = 7'h4c == auto_in_a_bits_source ? 5'h3 : _GEN_77; 
  assign _GEN_79 = 7'h4d == auto_in_a_bits_source ? 5'h3 : _GEN_78; 
  assign _GEN_80 = 7'h4e == auto_in_a_bits_source ? 5'h3 : _GEN_79; 
  assign _GEN_81 = 7'h4f == auto_in_a_bits_source ? 5'h3 : _GEN_80; 
  assign _GEN_82 = 7'h50 == auto_in_a_bits_source ? 5'h4 : _GEN_81; 
  assign _GEN_83 = 7'h51 == auto_in_a_bits_source ? 5'h4 : _GEN_82; 
  assign _GEN_84 = 7'h52 == auto_in_a_bits_source ? 5'h4 : _GEN_83; 
  assign _GEN_85 = 7'h53 == auto_in_a_bits_source ? 5'h4 : _GEN_84; 
  assign _GEN_86 = 7'h54 == auto_in_a_bits_source ? 5'h4 : _GEN_85; 
  assign _GEN_87 = 7'h55 == auto_in_a_bits_source ? 5'h4 : _GEN_86; 
  assign _GEN_88 = 7'h56 == auto_in_a_bits_source ? 5'h4 : _GEN_87; 
  assign _GEN_89 = 7'h57 == auto_in_a_bits_source ? 5'h4 : _GEN_88; 
  assign _GEN_90 = 7'h58 == auto_in_a_bits_source ? 5'h4 : _GEN_89; 
  assign _GEN_91 = 7'h59 == auto_in_a_bits_source ? 5'h4 : _GEN_90; 
  assign _GEN_92 = 7'h5a == auto_in_a_bits_source ? 5'h4 : _GEN_91; 
  assign _GEN_93 = 7'h5b == auto_in_a_bits_source ? 5'h4 : _GEN_92; 
  assign _GEN_94 = 7'h5c == auto_in_a_bits_source ? 5'h4 : _GEN_93; 
  assign _GEN_95 = 7'h5d == auto_in_a_bits_source ? 5'h4 : _GEN_94; 
  assign _GEN_96 = 7'h5e == auto_in_a_bits_source ? 5'h4 : _GEN_95; 
  assign _GEN_97 = 7'h5f == auto_in_a_bits_source ? 5'h4 : _GEN_96; 
  assign _GEN_98 = 7'h60 == auto_in_a_bits_source ? 5'h5 : _GEN_97; 
  assign _GEN_99 = 7'h61 == auto_in_a_bits_source ? 5'h5 : _GEN_98; 
  assign _GEN_100 = 7'h62 == auto_in_a_bits_source ? 5'h5 : _GEN_99; 
  assign _GEN_101 = 7'h63 == auto_in_a_bits_source ? 5'h5 : _GEN_100; 
  assign _GEN_102 = 7'h64 == auto_in_a_bits_source ? 5'h5 : _GEN_101; 
  assign _GEN_103 = 7'h65 == auto_in_a_bits_source ? 5'h5 : _GEN_102; 
  assign _GEN_104 = 7'h66 == auto_in_a_bits_source ? 5'h5 : _GEN_103; 
  assign _GEN_105 = 7'h67 == auto_in_a_bits_source ? 5'h5 : _GEN_104; 
  assign _GEN_106 = 7'h68 == auto_in_a_bits_source ? 5'h5 : _GEN_105; 
  assign _GEN_107 = 7'h69 == auto_in_a_bits_source ? 5'h5 : _GEN_106; 
  assign _GEN_108 = 7'h6a == auto_in_a_bits_source ? 5'h5 : _GEN_107; 
  assign _GEN_109 = 7'h6b == auto_in_a_bits_source ? 5'h5 : _GEN_108; 
  assign _GEN_110 = 7'h6c == auto_in_a_bits_source ? 5'h5 : _GEN_109; 
  assign _GEN_111 = 7'h6d == auto_in_a_bits_source ? 5'h5 : _GEN_110; 
  assign _GEN_112 = 7'h6e == auto_in_a_bits_source ? 5'h5 : _GEN_111; 
  assign _GEN_113 = 7'h6f == auto_in_a_bits_source ? 5'h5 : _GEN_112; 
  assign _GEN_114 = 7'h70 == auto_in_a_bits_source ? 5'h6 : _GEN_113; 
  assign _GEN_115 = 7'h71 == auto_in_a_bits_source ? 5'h6 : _GEN_114; 
  assign _GEN_116 = 7'h72 == auto_in_a_bits_source ? 5'h6 : _GEN_115; 
  assign _GEN_117 = 7'h73 == auto_in_a_bits_source ? 5'h6 : _GEN_116; 
  assign _GEN_118 = 7'h74 == auto_in_a_bits_source ? 5'h6 : _GEN_117; 
  assign _GEN_119 = 7'h75 == auto_in_a_bits_source ? 5'h6 : _GEN_118; 
  assign _GEN_120 = 7'h76 == auto_in_a_bits_source ? 5'h6 : _GEN_119; 
  assign _GEN_121 = 7'h77 == auto_in_a_bits_source ? 5'h6 : _GEN_120; 
  assign _GEN_122 = 7'h78 == auto_in_a_bits_source ? 5'h6 : _GEN_121; 
  assign _GEN_123 = 7'h79 == auto_in_a_bits_source ? 5'h6 : _GEN_122; 
  assign _GEN_124 = 7'h7a == auto_in_a_bits_source ? 5'h6 : _GEN_123; 
  assign _GEN_125 = 7'h7b == auto_in_a_bits_source ? 5'h6 : _GEN_124; 
  assign _GEN_126 = 7'h7c == auto_in_a_bits_source ? 5'h6 : _GEN_125; 
  assign _GEN_127 = 7'h7d == auto_in_a_bits_source ? 5'h6 : _GEN_126; 
  assign _GEN_128 = 7'h7e == auto_in_a_bits_source ? 5'h6 : _GEN_127; 
  assign _GEN_129 = 7'h7f == auto_in_a_bits_source ? 5'h6 : _GEN_128; 
  assign _T_61 = 18'h7ff << auto_in_a_bits_size; 
  assign _T_62 = _T_61[10:0]; 
  assign _T_63 = ~ _T_62; 
  assign _T_65 = auto_in_a_bits_size >= 3'h3; 
  assign _T_74 = _T_68 & auto_in_a_valid; 
  assign _T_75 = _T_57 == 1'h0; 
  assign _T_76 = _T_75 & _T_50_ready; 
  assign _T_77 = _T_13 ? _T_76 : 1'h1; 
  assign _T_78 = _T_74 & _T_77; 
  assign _T_81 = _T_74 & _T_13; 
  assign _T_85 = auto_in_d_ready & auto_out_rvalid; 
  assign _T_86 = auto_out_rlast == 1'h0; 
  assign _T_87 = auto_out_rvalid | _T_84; 
  assign _T_88 = _T_87 == 1'h0; 
  assign _T_90 = _T_87 ? auto_out_rvalid : auto_out_bvalid; 
  assign _T_93 = auto_out_rresp == 2'h3; 
  assign _GEN_260 = _T_91 ? _T_93 : _T_94; 
  assign _T_96 = auto_out_rresp != 2'h0; 
  assign _T_97 = auto_out_bresp != 2'h0; 
  assign _T_98 = _T_96 | _GEN_260; 
  assign _T_103 = 32'h1 << _GEN_129; 
  assign _T_104 = _T_103[22:0]; 
  assign _T_105 = _T_104[0]; 
  assign _T_106 = _T_104[1]; 
  assign _T_107 = _T_104[2]; 
  assign _T_108 = _T_104[3]; 
  assign _T_109 = _T_104[4]; 
  assign _T_110 = _T_104[5]; 
  assign _T_111 = _T_104[6]; 
  assign _T_112 = _T_104[7]; 
  assign _T_113 = _T_104[8]; 
  assign _T_114 = _T_104[9]; 
  assign _T_115 = _T_104[10]; 
  assign _T_116 = _T_104[11]; 
  assign _T_117 = _T_104[12]; 
  assign _T_118 = _T_104[13]; 
  assign _T_119 = _T_104[14]; 
  assign _T_120 = _T_104[15]; 
  assign _T_121 = _T_104[16]; 
  assign _T_122 = _T_104[17]; 
  assign _T_123 = _T_104[18]; 
  assign _T_124 = _T_104[19]; 
  assign _T_125 = _T_104[20]; 
  assign _T_126 = _T_104[21]; 
  assign _T_127 = _T_104[22]; 
  assign _T_128 = _T_87 ? auto_out_rid : auto_out_bid; 
  assign _T_130 = 32'h1 << _T_128; 
  assign _T_131 = _T_130[22:0]; 
  assign _T_132 = _T_131[0]; 
  assign _T_133 = _T_131[1]; 
  assign _T_134 = _T_131[2]; 
  assign _T_135 = _T_131[3]; 
  assign _T_136 = _T_131[4]; 
  assign _T_137 = _T_131[5]; 
  assign _T_138 = _T_131[6]; 
  assign _T_139 = _T_131[7]; 
  assign _T_140 = _T_131[8]; 
  assign _T_141 = _T_131[9]; 
  assign _T_142 = _T_131[10]; 
  assign _T_143 = _T_131[11]; 
  assign _T_144 = _T_131[12]; 
  assign _T_145 = _T_131[13]; 
  assign _T_146 = _T_131[14]; 
  assign _T_147 = _T_131[15]; 
  assign _T_148 = _T_131[16]; 
  assign _T_149 = _T_131[17]; 
  assign _T_150 = _T_131[18]; 
  assign _T_151 = _T_131[19]; 
  assign _T_152 = _T_131[20]; 
  assign _T_153 = _T_131[21]; 
  assign _T_154 = _T_131[22]; 
  assign _T_155 = _T_87 ? auto_out_rlast : 1'h1; 
  assign _T_159 = _T_49_ready & _T_78; 
  assign _T_160 = _T_105 & _T_159; 
  assign _T_161 = _T_132 & _T_155; 
  assign _T_162 = auto_in_d_ready & _T_90; 
  assign _T_163 = _T_161 & _T_162; 
  assign _GEN_285 = {{4'd0}, _T_160}; 
  assign _T_165 = _T_156 + _GEN_285; 
  assign _GEN_286 = {{4'd0}, _T_163}; 
  assign _T_167 = _T_165 - _GEN_286; 
  assign _T_168 = _T_163 == 1'h0; 
  assign _T_169 = _T_156 != 5'h0; 
  assign _T_170 = _T_168 | _T_169; 
  assign _T_172 = _T_170 | reset; 
  assign _T_173 = _T_172 == 1'h0; 
  assign _T_174 = _T_160 == 1'h0; 
  assign _T_175 = _T_156 != 5'h10; 
  assign _T_176 = _T_174 | _T_175; 
  assign _T_178 = _T_176 | reset; 
  assign _T_179 = _T_178 == 1'h0; 
  assign _T_189 = _T_106 & _T_159; 
  assign _T_190 = _T_133 & _T_155; 
  assign _T_192 = _T_190 & _T_162; 
  assign _GEN_287 = {{4'd0}, _T_189}; 
  assign _T_194 = _T_185 + _GEN_287; 
  assign _GEN_288 = {{4'd0}, _T_192}; 
  assign _T_196 = _T_194 - _GEN_288; 
  assign _T_197 = _T_192 == 1'h0; 
  assign _T_198 = _T_185 != 5'h0; 
  assign _T_199 = _T_197 | _T_198; 
  assign _T_201 = _T_199 | reset; 
  assign _T_202 = _T_201 == 1'h0; 
  assign _T_203 = _T_189 == 1'h0; 
  assign _T_204 = _T_185 != 5'h10; 
  assign _T_205 = _T_203 | _T_204; 
  assign _T_207 = _T_205 | reset; 
  assign _T_208 = _T_207 == 1'h0; 
  assign _T_218 = _T_107 & _T_159; 
  assign _T_219 = _T_134 & _T_155; 
  assign _T_221 = _T_219 & _T_162; 
  assign _GEN_289 = {{4'd0}, _T_218}; 
  assign _T_223 = _T_214 + _GEN_289; 
  assign _GEN_290 = {{4'd0}, _T_221}; 
  assign _T_225 = _T_223 - _GEN_290; 
  assign _T_226 = _T_221 == 1'h0; 
  assign _T_227 = _T_214 != 5'h0; 
  assign _T_228 = _T_226 | _T_227; 
  assign _T_230 = _T_228 | reset; 
  assign _T_231 = _T_230 == 1'h0; 
  assign _T_232 = _T_218 == 1'h0; 
  assign _T_233 = _T_214 != 5'h10; 
  assign _T_234 = _T_232 | _T_233; 
  assign _T_236 = _T_234 | reset; 
  assign _T_237 = _T_236 == 1'h0; 
  assign _T_247 = _T_108 & _T_159; 
  assign _T_248 = _T_135 & _T_155; 
  assign _T_250 = _T_248 & _T_162; 
  assign _GEN_291 = {{4'd0}, _T_247}; 
  assign _T_252 = _T_243 + _GEN_291; 
  assign _GEN_292 = {{4'd0}, _T_250}; 
  assign _T_254 = _T_252 - _GEN_292; 
  assign _T_255 = _T_250 == 1'h0; 
  assign _T_256 = _T_243 != 5'h0; 
  assign _T_257 = _T_255 | _T_256; 
  assign _T_259 = _T_257 | reset; 
  assign _T_260 = _T_259 == 1'h0; 
  assign _T_261 = _T_247 == 1'h0; 
  assign _T_262 = _T_243 != 5'h10; 
  assign _T_263 = _T_261 | _T_262; 
  assign _T_265 = _T_263 | reset; 
  assign _T_266 = _T_265 == 1'h0; 
  assign _T_276 = _T_109 & _T_159; 
  assign _T_277 = _T_136 & _T_155; 
  assign _T_279 = _T_277 & _T_162; 
  assign _GEN_293 = {{4'd0}, _T_276}; 
  assign _T_281 = _T_272 + _GEN_293; 
  assign _GEN_294 = {{4'd0}, _T_279}; 
  assign _T_283 = _T_281 - _GEN_294; 
  assign _T_284 = _T_279 == 1'h0; 
  assign _T_285 = _T_272 != 5'h0; 
  assign _T_286 = _T_284 | _T_285; 
  assign _T_288 = _T_286 | reset; 
  assign _T_289 = _T_288 == 1'h0; 
  assign _T_290 = _T_276 == 1'h0; 
  assign _T_291 = _T_272 != 5'h10; 
  assign _T_292 = _T_290 | _T_291; 
  assign _T_294 = _T_292 | reset; 
  assign _T_295 = _T_294 == 1'h0; 
  assign _T_305 = _T_110 & _T_159; 
  assign _T_306 = _T_137 & _T_155; 
  assign _T_308 = _T_306 & _T_162; 
  assign _GEN_295 = {{4'd0}, _T_305}; 
  assign _T_310 = _T_301 + _GEN_295; 
  assign _GEN_296 = {{4'd0}, _T_308}; 
  assign _T_312 = _T_310 - _GEN_296; 
  assign _T_313 = _T_308 == 1'h0; 
  assign _T_314 = _T_301 != 5'h0; 
  assign _T_315 = _T_313 | _T_314; 
  assign _T_317 = _T_315 | reset; 
  assign _T_318 = _T_317 == 1'h0; 
  assign _T_319 = _T_305 == 1'h0; 
  assign _T_320 = _T_301 != 5'h10; 
  assign _T_321 = _T_319 | _T_320; 
  assign _T_323 = _T_321 | reset; 
  assign _T_324 = _T_323 == 1'h0; 
  assign _T_334 = _T_111 & _T_159; 
  assign _T_335 = _T_138 & _T_155; 
  assign _T_337 = _T_335 & _T_162; 
  assign _GEN_297 = {{4'd0}, _T_334}; 
  assign _T_339 = _T_330 + _GEN_297; 
  assign _GEN_298 = {{4'd0}, _T_337}; 
  assign _T_341 = _T_339 - _GEN_298; 
  assign _T_342 = _T_337 == 1'h0; 
  assign _T_343 = _T_330 != 5'h0; 
  assign _T_344 = _T_342 | _T_343; 
  assign _T_346 = _T_344 | reset; 
  assign _T_347 = _T_346 == 1'h0; 
  assign _T_348 = _T_334 == 1'h0; 
  assign _T_349 = _T_330 != 5'h10; 
  assign _T_350 = _T_348 | _T_349; 
  assign _T_352 = _T_350 | reset; 
  assign _T_353 = _T_352 == 1'h0; 
  assign _T_363 = _T_112 & _T_159; 
  assign _T_364 = _T_139 & _T_155; 
  assign _T_366 = _T_364 & _T_162; 
  assign _T_368 = _T_359 + _T_363; 
  assign _T_370 = _T_368 - _T_366; 
  assign _T_371 = _T_366 == 1'h0; 
  assign _T_373 = _T_371 | _T_359; 
  assign _T_375 = _T_373 | reset; 
  assign _T_376 = _T_375 == 1'h0; 
  assign _T_377 = _T_363 == 1'h0; 
  assign _T_378 = _T_359 != 1'h1; 
  assign _T_379 = _T_377 | _T_378; 
  assign _T_381 = _T_379 | reset; 
  assign _T_382 = _T_381 == 1'h0; 
  assign _T_391 = _T_113 & _T_159; 
  assign _T_392 = _T_140 & _T_155; 
  assign _T_394 = _T_392 & _T_162; 
  assign _T_396 = _T_387 + _T_391; 
  assign _T_398 = _T_396 - _T_394; 
  assign _T_399 = _T_394 == 1'h0; 
  assign _T_401 = _T_399 | _T_387; 
  assign _T_403 = _T_401 | reset; 
  assign _T_404 = _T_403 == 1'h0; 
  assign _T_405 = _T_391 == 1'h0; 
  assign _T_406 = _T_387 != 1'h1; 
  assign _T_407 = _T_405 | _T_406; 
  assign _T_409 = _T_407 | reset; 
  assign _T_410 = _T_409 == 1'h0; 
  assign _T_419 = _T_114 & _T_159; 
  assign _T_420 = _T_141 & _T_155; 
  assign _T_422 = _T_420 & _T_162; 
  assign _T_424 = _T_415 + _T_419; 
  assign _T_426 = _T_424 - _T_422; 
  assign _T_427 = _T_422 == 1'h0; 
  assign _T_429 = _T_427 | _T_415; 
  assign _T_431 = _T_429 | reset; 
  assign _T_432 = _T_431 == 1'h0; 
  assign _T_433 = _T_419 == 1'h0; 
  assign _T_434 = _T_415 != 1'h1; 
  assign _T_435 = _T_433 | _T_434; 
  assign _T_437 = _T_435 | reset; 
  assign _T_438 = _T_437 == 1'h0; 
  assign _T_447 = _T_115 & _T_159; 
  assign _T_448 = _T_142 & _T_155; 
  assign _T_450 = _T_448 & _T_162; 
  assign _T_452 = _T_443 + _T_447; 
  assign _T_454 = _T_452 - _T_450; 
  assign _T_455 = _T_450 == 1'h0; 
  assign _T_457 = _T_455 | _T_443; 
  assign _T_459 = _T_457 | reset; 
  assign _T_460 = _T_459 == 1'h0; 
  assign _T_461 = _T_447 == 1'h0; 
  assign _T_462 = _T_443 != 1'h1; 
  assign _T_463 = _T_461 | _T_462; 
  assign _T_465 = _T_463 | reset; 
  assign _T_466 = _T_465 == 1'h0; 
  assign _T_475 = _T_116 & _T_159; 
  assign _T_476 = _T_143 & _T_155; 
  assign _T_478 = _T_476 & _T_162; 
  assign _T_480 = _T_471 + _T_475; 
  assign _T_482 = _T_480 - _T_478; 
  assign _T_483 = _T_478 == 1'h0; 
  assign _T_485 = _T_483 | _T_471; 
  assign _T_487 = _T_485 | reset; 
  assign _T_488 = _T_487 == 1'h0; 
  assign _T_489 = _T_475 == 1'h0; 
  assign _T_490 = _T_471 != 1'h1; 
  assign _T_491 = _T_489 | _T_490; 
  assign _T_493 = _T_491 | reset; 
  assign _T_494 = _T_493 == 1'h0; 
  assign _T_503 = _T_117 & _T_159; 
  assign _T_504 = _T_144 & _T_155; 
  assign _T_506 = _T_504 & _T_162; 
  assign _T_508 = _T_499 + _T_503; 
  assign _T_510 = _T_508 - _T_506; 
  assign _T_511 = _T_506 == 1'h0; 
  assign _T_513 = _T_511 | _T_499; 
  assign _T_515 = _T_513 | reset; 
  assign _T_516 = _T_515 == 1'h0; 
  assign _T_517 = _T_503 == 1'h0; 
  assign _T_518 = _T_499 != 1'h1; 
  assign _T_519 = _T_517 | _T_518; 
  assign _T_521 = _T_519 | reset; 
  assign _T_522 = _T_521 == 1'h0; 
  assign _T_531 = _T_118 & _T_159; 
  assign _T_532 = _T_145 & _T_155; 
  assign _T_534 = _T_532 & _T_162; 
  assign _T_536 = _T_527 + _T_531; 
  assign _T_538 = _T_536 - _T_534; 
  assign _T_539 = _T_534 == 1'h0; 
  assign _T_541 = _T_539 | _T_527; 
  assign _T_543 = _T_541 | reset; 
  assign _T_544 = _T_543 == 1'h0; 
  assign _T_545 = _T_531 == 1'h0; 
  assign _T_546 = _T_527 != 1'h1; 
  assign _T_547 = _T_545 | _T_546; 
  assign _T_549 = _T_547 | reset; 
  assign _T_550 = _T_549 == 1'h0; 
  assign _T_559 = _T_119 & _T_159; 
  assign _T_560 = _T_146 & _T_155; 
  assign _T_562 = _T_560 & _T_162; 
  assign _T_564 = _T_555 + _T_559; 
  assign _T_566 = _T_564 - _T_562; 
  assign _T_567 = _T_562 == 1'h0; 
  assign _T_569 = _T_567 | _T_555; 
  assign _T_571 = _T_569 | reset; 
  assign _T_572 = _T_571 == 1'h0; 
  assign _T_573 = _T_559 == 1'h0; 
  assign _T_574 = _T_555 != 1'h1; 
  assign _T_575 = _T_573 | _T_574; 
  assign _T_577 = _T_575 | reset; 
  assign _T_578 = _T_577 == 1'h0; 
  assign _T_587 = _T_120 & _T_159; 
  assign _T_588 = _T_147 & _T_155; 
  assign _T_590 = _T_588 & _T_162; 
  assign _T_592 = _T_583 + _T_587; 
  assign _T_594 = _T_592 - _T_590; 
  assign _T_595 = _T_590 == 1'h0; 
  assign _T_597 = _T_595 | _T_583; 
  assign _T_599 = _T_597 | reset; 
  assign _T_600 = _T_599 == 1'h0; 
  assign _T_601 = _T_587 == 1'h0; 
  assign _T_602 = _T_583 != 1'h1; 
  assign _T_603 = _T_601 | _T_602; 
  assign _T_605 = _T_603 | reset; 
  assign _T_606 = _T_605 == 1'h0; 
  assign _T_615 = _T_121 & _T_159; 
  assign _T_616 = _T_148 & _T_155; 
  assign _T_618 = _T_616 & _T_162; 
  assign _T_620 = _T_611 + _T_615; 
  assign _T_622 = _T_620 - _T_618; 
  assign _T_623 = _T_618 == 1'h0; 
  assign _T_625 = _T_623 | _T_611; 
  assign _T_627 = _T_625 | reset; 
  assign _T_628 = _T_627 == 1'h0; 
  assign _T_629 = _T_615 == 1'h0; 
  assign _T_630 = _T_611 != 1'h1; 
  assign _T_631 = _T_629 | _T_630; 
  assign _T_633 = _T_631 | reset; 
  assign _T_634 = _T_633 == 1'h0; 
  assign _T_643 = _T_122 & _T_159; 
  assign _T_644 = _T_149 & _T_155; 
  assign _T_646 = _T_644 & _T_162; 
  assign _T_648 = _T_639 + _T_643; 
  assign _T_650 = _T_648 - _T_646; 
  assign _T_651 = _T_646 == 1'h0; 
  assign _T_653 = _T_651 | _T_639; 
  assign _T_655 = _T_653 | reset; 
  assign _T_656 = _T_655 == 1'h0; 
  assign _T_657 = _T_643 == 1'h0; 
  assign _T_658 = _T_639 != 1'h1; 
  assign _T_659 = _T_657 | _T_658; 
  assign _T_661 = _T_659 | reset; 
  assign _T_662 = _T_661 == 1'h0; 
  assign _T_671 = _T_123 & _T_159; 
  assign _T_672 = _T_150 & _T_155; 
  assign _T_674 = _T_672 & _T_162; 
  assign _T_676 = _T_667 + _T_671; 
  assign _T_678 = _T_676 - _T_674; 
  assign _T_679 = _T_674 == 1'h0; 
  assign _T_681 = _T_679 | _T_667; 
  assign _T_683 = _T_681 | reset; 
  assign _T_684 = _T_683 == 1'h0; 
  assign _T_685 = _T_671 == 1'h0; 
  assign _T_686 = _T_667 != 1'h1; 
  assign _T_687 = _T_685 | _T_686; 
  assign _T_689 = _T_687 | reset; 
  assign _T_690 = _T_689 == 1'h0; 
  assign _T_699 = _T_124 & _T_159; 
  assign _T_700 = _T_151 & _T_155; 
  assign _T_702 = _T_700 & _T_162; 
  assign _T_704 = _T_695 + _T_699; 
  assign _T_706 = _T_704 - _T_702; 
  assign _T_707 = _T_702 == 1'h0; 
  assign _T_709 = _T_707 | _T_695; 
  assign _T_711 = _T_709 | reset; 
  assign _T_712 = _T_711 == 1'h0; 
  assign _T_713 = _T_699 == 1'h0; 
  assign _T_714 = _T_695 != 1'h1; 
  assign _T_715 = _T_713 | _T_714; 
  assign _T_717 = _T_715 | reset; 
  assign _T_718 = _T_717 == 1'h0; 
  assign _T_727 = _T_125 & _T_159; 
  assign _T_728 = _T_152 & _T_155; 
  assign _T_730 = _T_728 & _T_162; 
  assign _T_732 = _T_723 + _T_727; 
  assign _T_734 = _T_732 - _T_730; 
  assign _T_735 = _T_730 == 1'h0; 
  assign _T_737 = _T_735 | _T_723; 
  assign _T_739 = _T_737 | reset; 
  assign _T_740 = _T_739 == 1'h0; 
  assign _T_741 = _T_727 == 1'h0; 
  assign _T_742 = _T_723 != 1'h1; 
  assign _T_743 = _T_741 | _T_742; 
  assign _T_745 = _T_743 | reset; 
  assign _T_746 = _T_745 == 1'h0; 
  assign _T_755 = _T_126 & _T_159; 
  assign _T_756 = _T_153 & _T_155; 
  assign _T_758 = _T_756 & _T_162; 
  assign _T_760 = _T_751 + _T_755; 
  assign _T_762 = _T_760 - _T_758; 
  assign _T_763 = _T_758 == 1'h0; 
  assign _T_765 = _T_763 | _T_751; 
  assign _T_767 = _T_765 | reset; 
  assign _T_768 = _T_767 == 1'h0; 
  assign _T_769 = _T_755 == 1'h0; 
  assign _T_770 = _T_751 != 1'h1; 
  assign _T_771 = _T_769 | _T_770; 
  assign _T_773 = _T_771 | reset; 
  assign _T_774 = _T_773 == 1'h0; 
  assign _T_783 = _T_127 & _T_159; 
  assign _T_784 = _T_154 & _T_155; 
  assign _T_786 = _T_784 & _T_162; 
  assign _T_788 = _T_779 + _T_783; 
  assign _T_790 = _T_788 - _T_786; 
  assign _T_791 = _T_786 == 1'h0; 
  assign _T_793 = _T_791 | _T_779; 
  assign _T_795 = _T_793 | reset; 
  assign _T_796 = _T_795 == 1'h0; 
  assign _T_797 = _T_783 == 1'h0; 
  assign _T_798 = _T_779 != 1'h1; 
  assign _T_799 = _T_797 | _T_798; 
  assign _T_801 = _T_799 | reset; 
  assign _T_802 = _T_801 == 1'h0; 
  assign auto_in_a_ready = _T_68 & _T_71; 
  assign auto_in_d_valid = _T_87 ? auto_out_rvalid : auto_out_bvalid; 
  assign auto_in_d_bits_opcode = _T_87 ? 3'h1 : 3'h0; 
  assign auto_in_d_bits_size = _T_87 ? _T_46 : _T_48; 
  assign auto_in_d_bits_source = _T_87 ? _T_45 : _T_47; 
  assign auto_in_d_bits_denied = _T_87 ? _GEN_260 : _T_97; 
  assign auto_in_d_bits_data = auto_out_rdata; 
  assign auto_in_d_bits_corrupt = _T_87 ? _T_98 : 1'h0; 
  assign auto_out_awvalid = _T_52_valid & _T_52_bits_wen; 
  assign auto_out_awid = Queue_1_io_deq_bits_id; 
  assign auto_out_awaddr = Queue_1_io_deq_bits_addr; 
  assign auto_out_awlen = Queue_1_io_deq_bits_len; 
  assign auto_out_awsize = Queue_1_io_deq_bits_size; 
  assign auto_out_awburst = Queue_1_io_deq_bits_burst; 
  assign auto_out_awlock = Queue_1_io_deq_bits_lock; 
  assign auto_out_awcache = Queue_1_io_deq_bits_cache; 
  assign auto_out_awprot = Queue_1_io_deq_bits_prot; 
  assign auto_out_awqos = Queue_1_io_deq_bits_qos; 
  assign auto_out_awuser = Queue_1_io_deq_bits_user; 
  assign auto_out_awinstret = Queue_1_io_deq_bits_instret; 
  assign auto_out_wvalid = Queue_io_deq_valid; 
  assign auto_out_wdata = Queue_io_deq_bits_data; 
  assign auto_out_wstrb = Queue_io_deq_bits_strb; 
  assign auto_out_wlast = Queue_io_deq_bits_last; 
  assign auto_out_bready = auto_in_d_ready & _T_88; 
  assign auto_out_arvalid = _T_52_valid & _T_53; 
  assign auto_out_arid = Queue_1_io_deq_bits_id; 
  assign auto_out_araddr = Queue_1_io_deq_bits_addr; 
  assign auto_out_arlen = Queue_1_io_deq_bits_len; 
  assign auto_out_arsize = Queue_1_io_deq_bits_size; 
  assign auto_out_arburst = Queue_1_io_deq_bits_burst; 
  assign auto_out_arlock = Queue_1_io_deq_bits_lock; 
  assign auto_out_arcache = Queue_1_io_deq_bits_cache; 
  assign auto_out_arprot = Queue_1_io_deq_bits_prot; 
  assign auto_out_arqos = Queue_1_io_deq_bits_qos; 
  assign auto_out_aruser = Queue_1_io_deq_bits_user; 
  assign auto_out_arinstret = Queue_1_io_deq_bits_instret; 
  assign auto_out_rready = auto_in_d_ready; 
  assign TLMonitor_clock = clock; 
  assign TLMonitor_reset = reset; 
  assign TLMonitor_io_in_a_ready = _T_68 & _T_71; 
  assign TLMonitor_io_in_a_valid = auto_in_a_valid; 
  assign TLMonitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; 
  assign TLMonitor_io_in_a_bits_param = auto_in_a_bits_param; 
  assign TLMonitor_io_in_a_bits_size = auto_in_a_bits_size; 
  assign TLMonitor_io_in_a_bits_source = auto_in_a_bits_source; 
  assign TLMonitor_io_in_a_bits_address = auto_in_a_bits_address; 
  assign TLMonitor_io_in_a_bits_mask = auto_in_a_bits_mask; 
  assign TLMonitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; 
  assign TLMonitor_io_in_d_ready = auto_in_d_ready; 
  assign TLMonitor_io_in_d_valid = _T_87 ? auto_out_rvalid : auto_out_bvalid; 
  assign TLMonitor_io_in_d_bits_opcode = _T_87 ? 3'h1 : 3'h0; 
  assign TLMonitor_io_in_d_bits_size = _T_87 ? _T_46 : _T_48; 
  assign TLMonitor_io_in_d_bits_source = _T_87 ? _T_45 : _T_47; 
  assign TLMonitor_io_in_d_bits_denied = _T_87 ? _GEN_260 : _T_97; 
  assign TLMonitor_io_in_d_bits_corrupt = _T_87 ? _T_98 : 1'h0; 
  assign Queue_clock = clock; 
  assign Queue_reset = reset; 
  assign Queue_io_enq_valid = _T_81 & _T_69; 
  assign Queue_io_enq_bits_data = auto_in_a_bits_data; 
  assign Queue_io_enq_bits_strb = auto_in_a_bits_mask; 
  assign Queue_io_enq_bits_last = _T_27 | _T_28; 
  assign Queue_io_deq_ready = auto_out_wready; 
  assign Queue_1_clock = clock; 
  assign Queue_1_reset = reset; 
  assign Queue_1_io_enq_valid = _T_74 & _T_77; 
  assign Queue_1_io_enq_bits_id = 7'h7f == auto_in_a_bits_source ? 5'h6 : _GEN_128; 
  assign Queue_1_io_enq_bits_addr = auto_in_a_bits_address; 
  assign Queue_1_io_enq_bits_len = _T_63[10:3]; 
  assign Queue_1_io_enq_bits_size = _T_65 ? 3'h3 : auto_in_a_bits_size; 
  assign Queue_1_io_enq_bits_user = {{1'd0}, _T_44}; 
  assign Queue_1_io_enq_bits_wen = _T_12 == 1'h0; 
  assign Queue_1_io_deq_ready = _T_52_bits_wen ? auto_out_awready : auto_out_arready; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_330 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_331 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_301 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_302 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_272 = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_273 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_243 = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_244 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_214 = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_215 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_185 = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_186 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_156 = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_157 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_779 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_751 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_723 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_695 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_667 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_639 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_611 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_583 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_555 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_527 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_499 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_471 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_443 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_415 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_387 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_359 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_23 = _RAND_30[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_57 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_84 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_91 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_94 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_330 <= 5'h0;
    end else begin
      _T_330 <= _T_341;
    end
    if (_T_334) begin
      _T_331 <= _T_13;
    end
    if (reset) begin
      _T_301 <= 5'h0;
    end else begin
      _T_301 <= _T_312;
    end
    if (_T_305) begin
      _T_302 <= _T_13;
    end
    if (reset) begin
      _T_272 <= 5'h0;
    end else begin
      _T_272 <= _T_283;
    end
    if (_T_276) begin
      _T_273 <= _T_13;
    end
    if (reset) begin
      _T_243 <= 5'h0;
    end else begin
      _T_243 <= _T_254;
    end
    if (_T_247) begin
      _T_244 <= _T_13;
    end
    if (reset) begin
      _T_214 <= 5'h0;
    end else begin
      _T_214 <= _T_225;
    end
    if (_T_218) begin
      _T_215 <= _T_13;
    end
    if (reset) begin
      _T_185 <= 5'h0;
    end else begin
      _T_185 <= _T_196;
    end
    if (_T_189) begin
      _T_186 <= _T_13;
    end
    if (reset) begin
      _T_156 <= 5'h0;
    end else begin
      _T_156 <= _T_167;
    end
    if (_T_160) begin
      _T_157 <= _T_13;
    end
    if (reset) begin
      _T_779 <= 1'h0;
    end else begin
      _T_779 <= _T_790;
    end
    if (reset) begin
      _T_751 <= 1'h0;
    end else begin
      _T_751 <= _T_762;
    end
    if (reset) begin
      _T_723 <= 1'h0;
    end else begin
      _T_723 <= _T_734;
    end
    if (reset) begin
      _T_695 <= 1'h0;
    end else begin
      _T_695 <= _T_706;
    end
    if (reset) begin
      _T_667 <= 1'h0;
    end else begin
      _T_667 <= _T_678;
    end
    if (reset) begin
      _T_639 <= 1'h0;
    end else begin
      _T_639 <= _T_650;
    end
    if (reset) begin
      _T_611 <= 1'h0;
    end else begin
      _T_611 <= _T_622;
    end
    if (reset) begin
      _T_583 <= 1'h0;
    end else begin
      _T_583 <= _T_594;
    end
    if (reset) begin
      _T_555 <= 1'h0;
    end else begin
      _T_555 <= _T_566;
    end
    if (reset) begin
      _T_527 <= 1'h0;
    end else begin
      _T_527 <= _T_538;
    end
    if (reset) begin
      _T_499 <= 1'h0;
    end else begin
      _T_499 <= _T_510;
    end
    if (reset) begin
      _T_471 <= 1'h0;
    end else begin
      _T_471 <= _T_482;
    end
    if (reset) begin
      _T_443 <= 1'h0;
    end else begin
      _T_443 <= _T_454;
    end
    if (reset) begin
      _T_415 <= 1'h0;
    end else begin
      _T_415 <= _T_426;
    end
    if (reset) begin
      _T_387 <= 1'h0;
    end else begin
      _T_387 <= _T_398;
    end
    if (reset) begin
      _T_359 <= 1'h0;
    end else begin
      _T_359 <= _T_370;
    end
    if (reset) begin
      _T_23 <= 3'h0;
    end else begin
      if (_T_14) begin
        if (_T_26) begin
          if (_T_13) begin
            _T_23 <= _T_19;
          end else begin
            _T_23 <= 3'h0;
          end
        end else begin
          _T_23 <= _T_25;
        end
      end
    end
    if (reset) begin
      _T_57 <= 1'h0;
    end else begin
      if (_T_14) begin
        _T_57 <= _T_59;
      end
    end
    if (reset) begin
      _T_84 <= 1'h0;
    end else begin
      if (_T_85) begin
        _T_84 <= _T_86;
      end
    end
    if (reset) begin
      _T_91 <= 1'h1;
    end else begin
      if (_T_85) begin
        _T_91 <= auto_out_rlast;
      end
    end
    if (_T_91) begin
      _T_94 <= _T_93;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:125 assert (a_source  < UInt(BigInt(1) << sourceBits))\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:126 assert (a_size    < UInt(BigInt(1) << sizeBits))\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_173) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_173) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_179) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_179) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_202) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_202) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_208) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_208) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_231) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_231) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_237) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_237) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_260) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_260) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_266) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_266) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_289) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_289) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_295) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_295) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_318) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_318) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_324) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_324) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_347) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_347) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_353) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_353) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_376) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_376) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_382) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_382) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_404) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_404) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_410) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_410) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_432) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_432) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_438) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_438) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_460) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_460) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_466) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_466) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_488) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_488) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_494) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_494) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_516) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_516) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_522) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_522) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_544) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_544) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_550) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_550) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_572) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_572) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_578) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_578) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_600) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_600) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_606) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_606) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_628) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_628) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_634) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_634) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_656) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_656) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_662) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_662) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_684) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_684) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_690) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_690) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_712) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_712) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_718) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_718) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_740) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_740) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_746) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_746) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_768) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_768) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_774) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_774) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_796) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:233 assert (!dec || count =/= UInt(0))        // underflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_796) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_802) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:234 assert (!inc || count =/= UInt(maxCount)) // overflow\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_802) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLWidthWidget_1( 
  input         clock, 
  input         reset, 
  output        auto_in_a_ready, 
  input         auto_in_a_valid, 
  input  [2:0]  auto_in_a_bits_opcode, 
  input  [2:0]  auto_in_a_bits_param, 
  input  [3:0]  auto_in_a_bits_size, 
  input  [5:0]  auto_in_a_bits_source, 
  input  [31:0] auto_in_a_bits_address, 
  input  [3:0]  auto_in_a_bits_mask, 
  input  [31:0] auto_in_a_bits_data, 
  output        auto_in_c_ready, 
  input         auto_in_c_valid, 
  input  [2:0]  auto_in_c_bits_opcode, 
  input  [2:0]  auto_in_c_bits_param, 
  input  [3:0]  auto_in_c_bits_size, 
  input  [5:0]  auto_in_c_bits_source, 
  input  [31:0] auto_in_c_bits_address, 
  input         auto_in_c_bits_corrupt, 
  input         auto_in_d_ready, 
  output        auto_in_d_valid, 
  output [2:0]  auto_in_d_bits_opcode, 
  output [1:0]  auto_in_d_bits_param, 
  output [3:0]  auto_in_d_bits_size, 
  output [5:0]  auto_in_d_bits_source, 
  output        auto_in_d_bits_sink, 
  output        auto_in_d_bits_denied, 
  output [31:0] auto_in_d_bits_data, 
  output        auto_in_d_bits_corrupt, 
  output        auto_in_e_ready, 
  input         auto_in_e_valid, 
  input         auto_in_e_bits_sink, 
  input         auto_out_a_ready, 
  output        auto_out_a_valid, 
  output [2:0]  auto_out_a_bits_opcode, 
  output [2:0]  auto_out_a_bits_param, 
  output [3:0]  auto_out_a_bits_size, 
  output [5:0]  auto_out_a_bits_source, 
  output [31:0] auto_out_a_bits_address, 
  output [7:0]  auto_out_a_bits_mask, 
  output [63:0] auto_out_a_bits_data, 
  input         auto_out_c_ready, 
  output        auto_out_c_valid, 
  output [2:0]  auto_out_c_bits_opcode, 
  output [2:0]  auto_out_c_bits_param, 
  output [3:0]  auto_out_c_bits_size, 
  output [5:0]  auto_out_c_bits_source, 
  output [31:0] auto_out_c_bits_address, 
  output        auto_out_c_bits_corrupt, 
  output        auto_out_d_ready, 
  input         auto_out_d_valid, 
  input  [2:0]  auto_out_d_bits_opcode, 
  input  [1:0]  auto_out_d_bits_param, 
  input  [3:0]  auto_out_d_bits_size, 
  input  [5:0]  auto_out_d_bits_source, 
  input         auto_out_d_bits_sink, 
  input         auto_out_d_bits_denied, 
  input  [63:0] auto_out_d_bits_data, 
  input         auto_out_d_bits_corrupt, 
  input         auto_out_e_ready, 
  output        auto_out_e_valid, 
  output        auto_out_e_bits_sink 
);
  wire  TLMonitor_clock; 
  wire  TLMonitor_reset; 
  wire  TLMonitor_io_in_a_ready; 
  wire  TLMonitor_io_in_a_valid; 
  wire [2:0] TLMonitor_io_in_a_bits_opcode; 
  wire [2:0] TLMonitor_io_in_a_bits_param; 
  wire [3:0] TLMonitor_io_in_a_bits_size; 
  wire [5:0] TLMonitor_io_in_a_bits_source; 
  wire [31:0] TLMonitor_io_in_a_bits_address; 
  wire [3:0] TLMonitor_io_in_a_bits_mask; 
  wire  TLMonitor_io_in_c_ready; 
  wire  TLMonitor_io_in_c_valid; 
  wire [2:0] TLMonitor_io_in_c_bits_opcode; 
  wire [2:0] TLMonitor_io_in_c_bits_param; 
  wire [3:0] TLMonitor_io_in_c_bits_size; 
  wire [5:0] TLMonitor_io_in_c_bits_source; 
  wire [31:0] TLMonitor_io_in_c_bits_address; 
  wire  TLMonitor_io_in_c_bits_corrupt; 
  wire  TLMonitor_io_in_d_ready; 
  wire  TLMonitor_io_in_d_valid; 
  wire [2:0] TLMonitor_io_in_d_bits_opcode; 
  wire [1:0] TLMonitor_io_in_d_bits_param; 
  wire [3:0] TLMonitor_io_in_d_bits_size; 
  wire [5:0] TLMonitor_io_in_d_bits_source; 
  wire  TLMonitor_io_in_d_bits_sink; 
  wire  TLMonitor_io_in_d_bits_denied; 
  wire  TLMonitor_io_in_d_bits_corrupt; 
  wire  TLMonitor_io_in_e_ready; 
  wire  TLMonitor_io_in_e_valid; 
  wire  TLMonitor_io_in_e_bits_sink; 
  wire  Repeater_clock; 
  wire  Repeater_reset; 
  wire  Repeater_io_repeat; 
  wire  Repeater_io_enq_ready; 
  wire  Repeater_io_enq_valid; 
  wire [2:0] Repeater_io_enq_bits_opcode; 
  wire [1:0] Repeater_io_enq_bits_param; 
  wire [3:0] Repeater_io_enq_bits_size; 
  wire [5:0] Repeater_io_enq_bits_source; 
  wire  Repeater_io_enq_bits_sink; 
  wire  Repeater_io_enq_bits_denied; 
  wire [63:0] Repeater_io_enq_bits_data; 
  wire  Repeater_io_enq_bits_corrupt; 
  wire  Repeater_io_deq_ready; 
  wire  Repeater_io_deq_valid; 
  wire [2:0] Repeater_io_deq_bits_opcode; 
  wire [1:0] Repeater_io_deq_bits_param; 
  wire [3:0] Repeater_io_deq_bits_size; 
  wire [5:0] Repeater_io_deq_bits_source; 
  wire  Repeater_io_deq_bits_sink; 
  wire  Repeater_io_deq_bits_denied; 
  wire [63:0] Repeater_io_deq_bits_data; 
  wire  Repeater_io_deq_bits_corrupt; 
  wire  _T_8; 
  wire  _T_9; 
  wire [17:0] _T_11; 
  wire [2:0] _T_12; 
  wire [2:0] _T_13; 
  wire  _T_14; 
  reg  _T_15; 
  reg [31:0] _RAND_0;
  wire  _T_17; 
  wire  _T_18; 
  wire  _T_19; 
  wire  _T_21; 
  wire  _T_23; 
  wire  _T_33; 
  wire  _T_34; 
  wire  _T_30; 
  wire  _T_32; 
  reg [31:0] _T_36_0; 
  reg [31:0] _RAND_1;
  wire [31:0] _T_37; 
  wire  _T_41; 
  wire [1:0] _T_44; 
  wire [3:0] _T_45; 
  wire [2:0] _T_46; 
  wire [2:0] _T_47; 
  wire  _T_48; 
  wire  _T_49; 
  wire  _T_50; 
  wire  _T_51; 
  wire  _T_53; 
  wire  _T_54; 
  wire  _T_56; 
  wire  _T_57; 
  wire  _T_58; 
  wire  _T_59; 
  wire  _T_60; 
  wire  _T_61; 
  wire  _T_62; 
  wire  _T_63; 
  wire  _T_64; 
  wire  _T_65; 
  wire  _T_66; 
  wire  _T_67; 
  wire  _T_68; 
  wire  _T_69; 
  wire  _T_70; 
  wire  _T_71; 
  wire  _T_72; 
  wire  _T_73; 
  wire  _T_74; 
  wire  _T_75; 
  wire  _T_76; 
  wire  _T_77; 
  wire  _T_78; 
  wire  _T_79; 
  wire  _T_80; 
  wire  _T_81; 
  wire  _T_82; 
  wire  _T_83; 
  wire  _T_84; 
  wire  _T_85; 
  wire  _T_86; 
  wire  _T_87; 
  wire  _T_88; 
  wire  _T_89; 
  wire  _T_90; 
  wire  _T_91; 
  wire  _T_92; 
  wire  _T_93; 
  wire  _T_94; 
  wire  _T_95; 
  wire  _T_96; 
  wire  _T_97; 
  wire  _T_98; 
  wire  _T_99; 
  wire [7:0] _T_106; 
  reg [3:0] _T_107_0; 
  reg [31:0] _RAND_2;
  wire [3:0] _T_108; 
  wire [7:0] _T_113; 
  wire [7:0] _T_115; 
  wire [31:0] _T_119; 
  wire [31:0] _T_120; 
  wire [63:0] _T_121; 
  wire [2:0] _T_118_bits_opcode; 
  wire  _T_122; 
  wire [3:0] _T_118_bits_size; 
  wire [17:0] _T_124; 
  wire [2:0] _T_125; 
  wire [2:0] _T_126; 
  wire  _T_127; 
  reg  _T_128; 
  reg [31:0] _RAND_3;
  wire  _T_129; 
  wire  _T_130; 
  wire  _T_131; 
  wire  _T_132; 
  wire  _T_118_valid; 
  wire  _T_133; 
  wire  _T_135; 
  reg  _T_136_0; 
  reg [31:0] _RAND_4;
  reg  _T_136_1; 
  reg [31:0] _RAND_5;
  reg  _T_136_2; 
  reg [31:0] _RAND_6;
  reg  _T_136_3; 
  reg [31:0] _RAND_7;
  reg  _T_136_4; 
  reg [31:0] _RAND_8;
  reg  _T_136_5; 
  reg [31:0] _RAND_9;
  reg  _T_136_6; 
  reg [31:0] _RAND_10;
  reg  _T_136_7; 
  reg [31:0] _RAND_11;
  reg  _T_136_8; 
  reg [31:0] _RAND_12;
  reg  _T_136_9; 
  reg [31:0] _RAND_13;
  reg  _T_136_10; 
  reg [31:0] _RAND_14;
  reg  _T_136_11; 
  reg [31:0] _RAND_15;
  reg  _T_136_12; 
  reg [31:0] _RAND_16;
  reg  _T_136_13; 
  reg [31:0] _RAND_17;
  reg  _T_136_14; 
  reg [31:0] _RAND_18;
  reg  _T_136_15; 
  reg [31:0] _RAND_19;
  reg  _T_136_16; 
  reg [31:0] _RAND_20;
  reg  _T_136_17; 
  reg [31:0] _RAND_21;
  reg  _T_136_18; 
  reg [31:0] _RAND_22;
  reg  _T_136_19; 
  reg [31:0] _RAND_23;
  reg  _T_136_20; 
  reg [31:0] _RAND_24;
  reg  _T_136_21; 
  reg [31:0] _RAND_25;
  reg  _T_136_22; 
  reg [31:0] _RAND_26;
  reg  _T_136_23; 
  reg [31:0] _RAND_27;
  reg  _T_136_24; 
  reg [31:0] _RAND_28;
  reg  _T_136_25; 
  reg [31:0] _RAND_29;
  reg  _T_136_26; 
  reg [31:0] _RAND_30;
  reg  _T_136_27; 
  reg [31:0] _RAND_31;
  reg  _T_136_28; 
  reg [31:0] _RAND_32;
  reg  _T_136_29; 
  reg [31:0] _RAND_33;
  reg  _T_136_30; 
  reg [31:0] _RAND_34;
  reg  _T_136_31; 
  reg [31:0] _RAND_35;
  reg  _T_136_32; 
  reg [31:0] _RAND_36;
  reg  _T_136_33; 
  reg [31:0] _RAND_37;
  reg  _T_136_34; 
  reg [31:0] _RAND_38;
  reg  _T_136_35; 
  reg [31:0] _RAND_39;
  reg  _T_136_36; 
  reg [31:0] _RAND_40;
  reg  _T_136_37; 
  reg [31:0] _RAND_41;
  reg  _T_136_38; 
  reg [31:0] _RAND_42;
  reg  _T_136_39; 
  reg [31:0] _RAND_43;
  reg  _T_136_40; 
  reg [31:0] _RAND_44;
  reg  _T_136_41; 
  reg [31:0] _RAND_45;
  reg  _T_136_42; 
  reg [31:0] _RAND_46;
  reg  _T_136_43; 
  reg [31:0] _RAND_47;
  reg  _T_136_44; 
  reg [31:0] _RAND_48;
  reg  _T_136_45; 
  reg [31:0] _RAND_49;
  reg  _T_136_46; 
  reg [31:0] _RAND_50;
  reg  _T_136_47; 
  reg [31:0] _RAND_51;
  reg  _T_136_48; 
  reg [31:0] _RAND_52;
  reg  _T_136_49; 
  reg [31:0] _RAND_53;
  reg  _T_136_50; 
  reg [31:0] _RAND_54;
  reg  _T_136_51; 
  reg [31:0] _RAND_55;
  reg  _T_136_52; 
  reg [31:0] _RAND_56;
  reg  _T_136_53; 
  reg [31:0] _RAND_57;
  reg  _T_136_54; 
  reg [31:0] _RAND_58;
  reg  _T_136_55; 
  reg [31:0] _RAND_59;
  reg  _T_136_56; 
  reg [31:0] _RAND_60;
  reg  _T_136_57; 
  reg [31:0] _RAND_61;
  reg  _T_136_58; 
  reg [31:0] _RAND_62;
  reg  _T_136_59; 
  reg [31:0] _RAND_63;
  reg  _T_136_60; 
  reg [31:0] _RAND_64;
  reg  _T_136_61; 
  reg [31:0] _RAND_65;
  reg  _T_136_62; 
  reg [31:0] _RAND_66;
  reg  _T_136_63; 
  reg [31:0] _RAND_67;
  wire [5:0] _T_118_bits_source; 
  reg  _T_141; 
  reg [31:0] _RAND_68;
  wire  _GEN_137; 
  wire  _GEN_138; 
  wire  _GEN_139; 
  wire  _GEN_140; 
  wire  _GEN_141; 
  wire  _GEN_142; 
  wire  _GEN_143; 
  wire  _GEN_144; 
  wire  _GEN_145; 
  wire  _GEN_146; 
  wire  _GEN_147; 
  wire  _GEN_148; 
  wire  _GEN_149; 
  wire  _GEN_150; 
  wire  _GEN_151; 
  wire  _GEN_152; 
  wire  _GEN_153; 
  wire  _GEN_154; 
  wire  _GEN_155; 
  wire  _GEN_156; 
  wire  _GEN_157; 
  wire  _GEN_158; 
  wire  _GEN_159; 
  wire  _GEN_160; 
  wire  _GEN_161; 
  wire  _GEN_162; 
  wire  _GEN_163; 
  wire  _GEN_164; 
  wire  _GEN_165; 
  wire  _GEN_166; 
  wire  _GEN_167; 
  wire  _GEN_168; 
  wire  _GEN_169; 
  wire  _GEN_170; 
  wire  _GEN_171; 
  wire  _GEN_172; 
  wire  _GEN_173; 
  wire  _GEN_174; 
  wire  _GEN_175; 
  wire  _GEN_176; 
  wire  _GEN_177; 
  wire  _GEN_178; 
  wire  _GEN_179; 
  wire  _GEN_180; 
  wire  _GEN_181; 
  wire  _GEN_182; 
  wire  _GEN_183; 
  wire  _GEN_184; 
  wire  _GEN_185; 
  wire  _GEN_186; 
  wire  _GEN_187; 
  wire  _GEN_188; 
  wire  _GEN_189; 
  wire  _GEN_190; 
  wire  _GEN_191; 
  wire  _GEN_192; 
  wire  _GEN_193; 
  wire  _GEN_194; 
  wire  _GEN_195; 
  wire  _GEN_196; 
  wire  _GEN_197; 
  wire  _GEN_198; 
  wire  _GEN_199; 
  wire  _GEN_200; 
  wire  _T_143; 
  wire  _T_144; 
  wire  _T_145; 
  wire [31:0] _T_146; 
  wire [31:0] _T_147; 
  wire  _T_176; 
  wire [17:0] _T_178; 
  wire [2:0] _T_179; 
  wire [2:0] _T_180; 
  wire  _T_181; 
  reg  _T_182; 
  reg [31:0] _RAND_69;
  wire  _T_184; 
  wire  _T_185; 
  wire  _T_186; 
  reg  _T_195; 
  reg [31:0] _RAND_70;
  wire  _T_196; 
  wire  _T_200; 
  wire  _T_201; 
  wire  _T_197; 
  wire  _T_199; 
  dual_TLMonitor_17 dual_TLMonitor ( 
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_c_ready(TLMonitor_io_in_c_ready),
    .io_in_c_valid(TLMonitor_io_in_c_valid),
    .io_in_c_bits_opcode(TLMonitor_io_in_c_bits_opcode),
    .io_in_c_bits_param(TLMonitor_io_in_c_bits_param),
    .io_in_c_bits_size(TLMonitor_io_in_c_bits_size),
    .io_in_c_bits_source(TLMonitor_io_in_c_bits_source),
    .io_in_c_bits_address(TLMonitor_io_in_c_bits_address),
    .io_in_c_bits_corrupt(TLMonitor_io_in_c_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt),
    .io_in_e_ready(TLMonitor_io_in_e_ready),
    .io_in_e_valid(TLMonitor_io_in_e_valid),
    .io_in_e_bits_sink(TLMonitor_io_in_e_bits_sink)
  );
  dual_Repeater_2 dual_Repeater_top ( 
    .clock(Repeater_clock),
    .reset(Repeater_reset),
    .io_repeat(Repeater_io_repeat),
    .io_enq_ready(Repeater_io_enq_ready),
    .io_enq_valid(Repeater_io_enq_valid),
    .io_enq_bits_opcode(Repeater_io_enq_bits_opcode),
    .io_enq_bits_param(Repeater_io_enq_bits_param),
    .io_enq_bits_size(Repeater_io_enq_bits_size),
    .io_enq_bits_source(Repeater_io_enq_bits_source),
    .io_enq_bits_sink(Repeater_io_enq_bits_sink),
    .io_enq_bits_denied(Repeater_io_enq_bits_denied),
    .io_enq_bits_data(Repeater_io_enq_bits_data),
    .io_enq_bits_corrupt(Repeater_io_enq_bits_corrupt),
    .io_deq_ready(Repeater_io_deq_ready),
    .io_deq_valid(Repeater_io_deq_valid),
    .io_deq_bits_opcode(Repeater_io_deq_bits_opcode),
    .io_deq_bits_param(Repeater_io_deq_bits_param),
    .io_deq_bits_size(Repeater_io_deq_bits_size),
    .io_deq_bits_source(Repeater_io_deq_bits_source),
    .io_deq_bits_sink(Repeater_io_deq_bits_sink),
    .io_deq_bits_denied(Repeater_io_deq_bits_denied),
    .io_deq_bits_data(Repeater_io_deq_bits_data),
    .io_deq_bits_corrupt(Repeater_io_deq_bits_corrupt)
  );
  assign _T_8 = auto_in_a_bits_opcode[2]; 
  assign _T_9 = _T_8 == 1'h0; 
  assign _T_11 = 18'h7 << auto_in_a_bits_size; 
  assign _T_12 = _T_11[2:0]; 
  assign _T_13 = ~ _T_12; 
  assign _T_14 = _T_13[2:2]; 
  assign _T_17 = _T_15 == _T_14; 
  assign _T_18 = _T_9 == 1'h0; 
  assign _T_19 = _T_17 | _T_18; 
  assign _T_21 = _T_15 & _T_14; 
  assign _T_23 = _T_21 == 1'h0; 
  assign _T_33 = _T_19 == 1'h0; 
  assign _T_34 = auto_out_a_ready | _T_33; 
  assign _T_30 = _T_34 & auto_in_a_valid; 
  assign _T_32 = _T_15 + 1'h1; 
  assign _T_37 = _T_23 ? auto_in_a_bits_data : _T_36_0; 
  assign _T_41 = _T_30 & _T_33; 
  assign _T_44 = auto_in_a_bits_size[1:0]; 
  assign _T_45 = 4'h1 << _T_44; 
  assign _T_46 = _T_45[2:0]; 
  assign _T_47 = _T_46 | 3'h1; 
  assign _T_48 = auto_in_a_bits_size >= 4'h3; 
  assign _T_49 = _T_47[2]; 
  assign _T_50 = auto_in_a_bits_address[2]; 
  assign _T_51 = _T_50 == 1'h0; 
  assign _T_53 = _T_49 & _T_51; 
  assign _T_54 = _T_48 | _T_53; 
  assign _T_56 = _T_49 & _T_50; 
  assign _T_57 = _T_48 | _T_56; 
  assign _T_58 = _T_47[1]; 
  assign _T_59 = auto_in_a_bits_address[1]; 
  assign _T_60 = _T_59 == 1'h0; 
  assign _T_61 = _T_51 & _T_60; 
  assign _T_62 = _T_58 & _T_61; 
  assign _T_63 = _T_54 | _T_62; 
  assign _T_64 = _T_51 & _T_59; 
  assign _T_65 = _T_58 & _T_64; 
  assign _T_66 = _T_54 | _T_65; 
  assign _T_67 = _T_50 & _T_60; 
  assign _T_68 = _T_58 & _T_67; 
  assign _T_69 = _T_57 | _T_68; 
  assign _T_70 = _T_50 & _T_59; 
  assign _T_71 = _T_58 & _T_70; 
  assign _T_72 = _T_57 | _T_71; 
  assign _T_73 = _T_47[0]; 
  assign _T_74 = auto_in_a_bits_address[0]; 
  assign _T_75 = _T_74 == 1'h0; 
  assign _T_76 = _T_61 & _T_75; 
  assign _T_77 = _T_73 & _T_76; 
  assign _T_78 = _T_63 | _T_77; 
  assign _T_79 = _T_61 & _T_74; 
  assign _T_80 = _T_73 & _T_79; 
  assign _T_81 = _T_63 | _T_80; 
  assign _T_82 = _T_64 & _T_75; 
  assign _T_83 = _T_73 & _T_82; 
  assign _T_84 = _T_66 | _T_83; 
  assign _T_85 = _T_64 & _T_74; 
  assign _T_86 = _T_73 & _T_85; 
  assign _T_87 = _T_66 | _T_86; 
  assign _T_88 = _T_67 & _T_75; 
  assign _T_89 = _T_73 & _T_88; 
  assign _T_90 = _T_69 | _T_89; 
  assign _T_91 = _T_67 & _T_74; 
  assign _T_92 = _T_73 & _T_91; 
  assign _T_93 = _T_69 | _T_92; 
  assign _T_94 = _T_70 & _T_75; 
  assign _T_95 = _T_73 & _T_94; 
  assign _T_96 = _T_72 | _T_95; 
  assign _T_97 = _T_70 & _T_74; 
  assign _T_98 = _T_73 & _T_97; 
  assign _T_99 = _T_72 | _T_98; 
  assign _T_106 = {_T_99,_T_96,_T_93,_T_90,_T_87,_T_84,_T_81,_T_78}; 
  assign _T_108 = _T_23 ? auto_in_a_bits_mask : _T_107_0; 
  assign _T_113 = {auto_in_a_bits_mask,_T_108}; 
  assign _T_115 = _T_9 ? _T_113 : 8'hff; 
  assign _T_119 = Repeater_io_deq_bits_data[63:32]; 
  assign _T_120 = auto_out_d_bits_data[31:0]; 
  assign _T_121 = {_T_119,_T_120}; 
  assign _T_118_bits_opcode = Repeater_io_deq_bits_opcode; 
  assign _T_122 = _T_118_bits_opcode[0]; 
  assign _T_118_bits_size = Repeater_io_deq_bits_size; 
  assign _T_124 = 18'h7 << _T_118_bits_size; 
  assign _T_125 = _T_124[2:0]; 
  assign _T_126 = ~ _T_125; 
  assign _T_127 = _T_126[2:2]; 
  assign _T_129 = _T_128 == 1'h0; 
  assign _T_130 = _T_128 == _T_127; 
  assign _T_131 = _T_122 == 1'h0; 
  assign _T_132 = _T_130 | _T_131; 
  assign _T_118_valid = Repeater_io_deq_valid; 
  assign _T_133 = auto_in_d_ready & _T_118_valid; 
  assign _T_135 = _T_128 + 1'h1; 
  assign _T_118_bits_source = Repeater_io_deq_bits_source; 
  assign _GEN_137 = 6'h1 == _T_118_bits_source ? _T_136_1 : _T_136_0; 
  assign _GEN_138 = 6'h2 == _T_118_bits_source ? _T_136_2 : _GEN_137; 
  assign _GEN_139 = 6'h3 == _T_118_bits_source ? _T_136_3 : _GEN_138; 
  assign _GEN_140 = 6'h4 == _T_118_bits_source ? _T_136_4 : _GEN_139; 
  assign _GEN_141 = 6'h5 == _T_118_bits_source ? _T_136_5 : _GEN_140; 
  assign _GEN_142 = 6'h6 == _T_118_bits_source ? _T_136_6 : _GEN_141; 
  assign _GEN_143 = 6'h7 == _T_118_bits_source ? _T_136_7 : _GEN_142; 
  assign _GEN_144 = 6'h8 == _T_118_bits_source ? _T_136_8 : _GEN_143; 
  assign _GEN_145 = 6'h9 == _T_118_bits_source ? _T_136_9 : _GEN_144; 
  assign _GEN_146 = 6'ha == _T_118_bits_source ? _T_136_10 : _GEN_145; 
  assign _GEN_147 = 6'hb == _T_118_bits_source ? _T_136_11 : _GEN_146; 
  assign _GEN_148 = 6'hc == _T_118_bits_source ? _T_136_12 : _GEN_147; 
  assign _GEN_149 = 6'hd == _T_118_bits_source ? _T_136_13 : _GEN_148; 
  assign _GEN_150 = 6'he == _T_118_bits_source ? _T_136_14 : _GEN_149; 
  assign _GEN_151 = 6'hf == _T_118_bits_source ? _T_136_15 : _GEN_150; 
  assign _GEN_152 = 6'h10 == _T_118_bits_source ? _T_136_16 : _GEN_151; 
  assign _GEN_153 = 6'h11 == _T_118_bits_source ? _T_136_17 : _GEN_152; 
  assign _GEN_154 = 6'h12 == _T_118_bits_source ? _T_136_18 : _GEN_153; 
  assign _GEN_155 = 6'h13 == _T_118_bits_source ? _T_136_19 : _GEN_154; 
  assign _GEN_156 = 6'h14 == _T_118_bits_source ? _T_136_20 : _GEN_155; 
  assign _GEN_157 = 6'h15 == _T_118_bits_source ? _T_136_21 : _GEN_156; 
  assign _GEN_158 = 6'h16 == _T_118_bits_source ? _T_136_22 : _GEN_157; 
  assign _GEN_159 = 6'h17 == _T_118_bits_source ? _T_136_23 : _GEN_158; 
  assign _GEN_160 = 6'h18 == _T_118_bits_source ? _T_136_24 : _GEN_159; 
  assign _GEN_161 = 6'h19 == _T_118_bits_source ? _T_136_25 : _GEN_160; 
  assign _GEN_162 = 6'h1a == _T_118_bits_source ? _T_136_26 : _GEN_161; 
  assign _GEN_163 = 6'h1b == _T_118_bits_source ? _T_136_27 : _GEN_162; 
  assign _GEN_164 = 6'h1c == _T_118_bits_source ? _T_136_28 : _GEN_163; 
  assign _GEN_165 = 6'h1d == _T_118_bits_source ? _T_136_29 : _GEN_164; 
  assign _GEN_166 = 6'h1e == _T_118_bits_source ? _T_136_30 : _GEN_165; 
  assign _GEN_167 = 6'h1f == _T_118_bits_source ? _T_136_31 : _GEN_166; 
  assign _GEN_168 = 6'h20 == _T_118_bits_source ? _T_136_32 : _GEN_167; 
  assign _GEN_169 = 6'h21 == _T_118_bits_source ? _T_136_33 : _GEN_168; 
  assign _GEN_170 = 6'h22 == _T_118_bits_source ? _T_136_34 : _GEN_169; 
  assign _GEN_171 = 6'h23 == _T_118_bits_source ? _T_136_35 : _GEN_170; 
  assign _GEN_172 = 6'h24 == _T_118_bits_source ? _T_136_36 : _GEN_171; 
  assign _GEN_173 = 6'h25 == _T_118_bits_source ? _T_136_37 : _GEN_172; 
  assign _GEN_174 = 6'h26 == _T_118_bits_source ? _T_136_38 : _GEN_173; 
  assign _GEN_175 = 6'h27 == _T_118_bits_source ? _T_136_39 : _GEN_174; 
  assign _GEN_176 = 6'h28 == _T_118_bits_source ? _T_136_40 : _GEN_175; 
  assign _GEN_177 = 6'h29 == _T_118_bits_source ? _T_136_41 : _GEN_176; 
  assign _GEN_178 = 6'h2a == _T_118_bits_source ? _T_136_42 : _GEN_177; 
  assign _GEN_179 = 6'h2b == _T_118_bits_source ? _T_136_43 : _GEN_178; 
  assign _GEN_180 = 6'h2c == _T_118_bits_source ? _T_136_44 : _GEN_179; 
  assign _GEN_181 = 6'h2d == _T_118_bits_source ? _T_136_45 : _GEN_180; 
  assign _GEN_182 = 6'h2e == _T_118_bits_source ? _T_136_46 : _GEN_181; 
  assign _GEN_183 = 6'h2f == _T_118_bits_source ? _T_136_47 : _GEN_182; 
  assign _GEN_184 = 6'h30 == _T_118_bits_source ? _T_136_48 : _GEN_183; 
  assign _GEN_185 = 6'h31 == _T_118_bits_source ? _T_136_49 : _GEN_184; 
  assign _GEN_186 = 6'h32 == _T_118_bits_source ? _T_136_50 : _GEN_185; 
  assign _GEN_187 = 6'h33 == _T_118_bits_source ? _T_136_51 : _GEN_186; 
  assign _GEN_188 = 6'h34 == _T_118_bits_source ? _T_136_52 : _GEN_187; 
  assign _GEN_189 = 6'h35 == _T_118_bits_source ? _T_136_53 : _GEN_188; 
  assign _GEN_190 = 6'h36 == _T_118_bits_source ? _T_136_54 : _GEN_189; 
  assign _GEN_191 = 6'h37 == _T_118_bits_source ? _T_136_55 : _GEN_190; 
  assign _GEN_192 = 6'h38 == _T_118_bits_source ? _T_136_56 : _GEN_191; 
  assign _GEN_193 = 6'h39 == _T_118_bits_source ? _T_136_57 : _GEN_192; 
  assign _GEN_194 = 6'h3a == _T_118_bits_source ? _T_136_58 : _GEN_193; 
  assign _GEN_195 = 6'h3b == _T_118_bits_source ? _T_136_59 : _GEN_194; 
  assign _GEN_196 = 6'h3c == _T_118_bits_source ? _T_136_60 : _GEN_195; 
  assign _GEN_197 = 6'h3d == _T_118_bits_source ? _T_136_61 : _GEN_196; 
  assign _GEN_198 = 6'h3e == _T_118_bits_source ? _T_136_62 : _GEN_197; 
  assign _GEN_199 = 6'h3f == _T_118_bits_source ? _T_136_63 : _GEN_198; 
  assign _GEN_200 = _T_129 ? _GEN_199 : _T_141; 
  assign _T_143 = ~ _T_127; 
  assign _T_144 = _GEN_200 & _T_143; 
  assign _T_145 = _T_144 | _T_128; 
  assign _T_146 = _T_121[31:0]; 
  assign _T_147 = _T_121[63:32]; 
  assign _T_176 = auto_in_c_bits_opcode[0]; 
  assign _T_178 = 18'h7 << auto_in_c_bits_size; 
  assign _T_179 = _T_178[2:0]; 
  assign _T_180 = ~ _T_179; 
  assign _T_181 = _T_180[2:2]; 
  assign _T_184 = _T_182 == _T_181; 
  assign _T_185 = _T_176 == 1'h0; 
  assign _T_186 = _T_184 | _T_185; 
  assign _T_196 = auto_in_c_bits_corrupt | _T_195; 
  assign _T_200 = _T_186 == 1'h0; 
  assign _T_201 = auto_out_c_ready | _T_200; 
  assign _T_197 = _T_201 & auto_in_c_valid; 
  assign _T_199 = _T_182 + 1'h1; 
  assign auto_in_a_ready = auto_out_a_ready | _T_33; 
  assign auto_in_c_ready = auto_out_c_ready | _T_200; 
  assign auto_in_d_valid = Repeater_io_deq_valid; 
  assign auto_in_d_bits_opcode = Repeater_io_deq_bits_opcode; 
  assign auto_in_d_bits_param = Repeater_io_deq_bits_param; 
  assign auto_in_d_bits_size = Repeater_io_deq_bits_size; 
  assign auto_in_d_bits_source = Repeater_io_deq_bits_source; 
  assign auto_in_d_bits_sink = Repeater_io_deq_bits_sink; 
  assign auto_in_d_bits_denied = Repeater_io_deq_bits_denied; 
  assign auto_in_d_bits_data = _T_145 ? _T_147 : _T_146; 
  assign auto_in_d_bits_corrupt = Repeater_io_deq_bits_corrupt; 
  assign auto_in_e_ready = auto_out_e_ready; 
  assign auto_out_a_valid = auto_in_a_valid & _T_19; 
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; 
  assign auto_out_a_bits_param = auto_in_a_bits_param; 
  assign auto_out_a_bits_size = auto_in_a_bits_size; 
  assign auto_out_a_bits_source = auto_in_a_bits_source; 
  assign auto_out_a_bits_address = auto_in_a_bits_address; 
  assign auto_out_a_bits_mask = _T_106 & _T_115; 
  assign auto_out_a_bits_data = {auto_in_a_bits_data,_T_37}; 
  assign auto_out_c_valid = auto_in_c_valid & _T_186; 
  assign auto_out_c_bits_opcode = auto_in_c_bits_opcode; 
  assign auto_out_c_bits_param = auto_in_c_bits_param; 
  assign auto_out_c_bits_size = auto_in_c_bits_size; 
  assign auto_out_c_bits_source = auto_in_c_bits_source; 
  assign auto_out_c_bits_address = auto_in_c_bits_address; 
  assign auto_out_c_bits_corrupt = auto_in_c_bits_corrupt | _T_195; 
  assign auto_out_d_ready = Repeater_io_enq_ready; 
  assign auto_out_e_valid = auto_in_e_valid; 
  assign auto_out_e_bits_sink = auto_in_e_bits_sink; 
  assign TLMonitor_clock = clock; 
  assign TLMonitor_reset = reset; 
  assign TLMonitor_io_in_a_ready = auto_out_a_ready | _T_33; 
  assign TLMonitor_io_in_a_valid = auto_in_a_valid; 
  assign TLMonitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; 
  assign TLMonitor_io_in_a_bits_param = auto_in_a_bits_param; 
  assign TLMonitor_io_in_a_bits_size = auto_in_a_bits_size; 
  assign TLMonitor_io_in_a_bits_source = auto_in_a_bits_source; 
  assign TLMonitor_io_in_a_bits_address = auto_in_a_bits_address; 
  assign TLMonitor_io_in_a_bits_mask = auto_in_a_bits_mask; 
  assign TLMonitor_io_in_c_ready = auto_out_c_ready | _T_200; 
  assign TLMonitor_io_in_c_valid = auto_in_c_valid; 
  assign TLMonitor_io_in_c_bits_opcode = auto_in_c_bits_opcode; 
  assign TLMonitor_io_in_c_bits_param = auto_in_c_bits_param; 
  assign TLMonitor_io_in_c_bits_size = auto_in_c_bits_size; 
  assign TLMonitor_io_in_c_bits_source = auto_in_c_bits_source; 
  assign TLMonitor_io_in_c_bits_address = auto_in_c_bits_address; 
  assign TLMonitor_io_in_c_bits_corrupt = auto_in_c_bits_corrupt; 
  assign TLMonitor_io_in_d_ready = auto_in_d_ready; 
  assign TLMonitor_io_in_d_valid = Repeater_io_deq_valid; 
  assign TLMonitor_io_in_d_bits_opcode = Repeater_io_deq_bits_opcode; 
  assign TLMonitor_io_in_d_bits_param = Repeater_io_deq_bits_param; 
  assign TLMonitor_io_in_d_bits_size = Repeater_io_deq_bits_size; 
  assign TLMonitor_io_in_d_bits_source = Repeater_io_deq_bits_source; 
  assign TLMonitor_io_in_d_bits_sink = Repeater_io_deq_bits_sink; 
  assign TLMonitor_io_in_d_bits_denied = Repeater_io_deq_bits_denied; 
  assign TLMonitor_io_in_d_bits_corrupt = Repeater_io_deq_bits_corrupt; 
  assign TLMonitor_io_in_e_ready = auto_out_e_ready; 
  assign TLMonitor_io_in_e_valid = auto_in_e_valid; 
  assign TLMonitor_io_in_e_bits_sink = auto_in_e_bits_sink; 
  assign Repeater_clock = clock; 
  assign Repeater_reset = reset; 
  assign Repeater_io_repeat = _T_132 == 1'h0; 
  assign Repeater_io_enq_valid = auto_out_d_valid; 
  assign Repeater_io_enq_bits_opcode = auto_out_d_bits_opcode; 
  assign Repeater_io_enq_bits_param = auto_out_d_bits_param; 
  assign Repeater_io_enq_bits_size = auto_out_d_bits_size; 
  assign Repeater_io_enq_bits_source = auto_out_d_bits_source; 
  assign Repeater_io_enq_bits_sink = auto_out_d_bits_sink; 
  assign Repeater_io_enq_bits_denied = auto_out_d_bits_denied; 
  assign Repeater_io_enq_bits_data = auto_out_d_bits_data; 
  assign Repeater_io_enq_bits_corrupt = auto_out_d_bits_corrupt; 
  assign Repeater_io_deq_ready = auto_in_d_ready; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_36_0 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_107_0 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_128 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_136_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_136_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_136_2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_136_3 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_136_4 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_136_5 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_136_6 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_136_7 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_136_8 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_136_9 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_136_10 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_136_11 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_136_12 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_136_13 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_136_14 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_136_15 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_136_16 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_136_17 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_136_18 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_136_19 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_136_20 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_136_21 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_136_22 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_136_23 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_136_24 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_136_25 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_136_26 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_136_27 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_136_28 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_136_29 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_136_30 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_136_31 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_136_32 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_136_33 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_136_34 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_136_35 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_136_36 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_136_37 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_136_38 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_136_39 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_136_40 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_136_41 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_136_42 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_136_43 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_136_44 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_136_45 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_136_46 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_136_47 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_136_48 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_136_49 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_136_50 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_136_51 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_136_52 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_136_53 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_136_54 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_136_55 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_136_56 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_136_57 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_136_58 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_136_59 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_136_60 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_136_61 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_136_62 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_136_63 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_141 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_182 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_195 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (_T_30) begin
        if (_T_19) begin
          _T_15 <= 1'h0;
        end else begin
          _T_15 <= _T_32;
        end
      end
    end
    if (_T_41) begin
      if (_T_23) begin
        _T_36_0 <= auto_in_a_bits_data;
      end
    end
    if (_T_41) begin
      if (_T_23) begin
        _T_107_0 <= auto_in_a_bits_mask;
      end
    end
    if (reset) begin
      _T_128 <= 1'h0;
    end else begin
      if (_T_133) begin
        if (_T_132) begin
          _T_128 <= 1'h0;
        end else begin
          _T_128 <= _T_135;
        end
      end
    end
    if (_T_30) begin
      if (6'h0 == auto_in_a_bits_source) begin
        _T_136_0 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h1 == auto_in_a_bits_source) begin
        _T_136_1 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h2 == auto_in_a_bits_source) begin
        _T_136_2 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h3 == auto_in_a_bits_source) begin
        _T_136_3 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h4 == auto_in_a_bits_source) begin
        _T_136_4 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h5 == auto_in_a_bits_source) begin
        _T_136_5 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h6 == auto_in_a_bits_source) begin
        _T_136_6 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h7 == auto_in_a_bits_source) begin
        _T_136_7 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h8 == auto_in_a_bits_source) begin
        _T_136_8 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h9 == auto_in_a_bits_source) begin
        _T_136_9 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'ha == auto_in_a_bits_source) begin
        _T_136_10 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'hb == auto_in_a_bits_source) begin
        _T_136_11 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'hc == auto_in_a_bits_source) begin
        _T_136_12 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'hd == auto_in_a_bits_source) begin
        _T_136_13 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'he == auto_in_a_bits_source) begin
        _T_136_14 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'hf == auto_in_a_bits_source) begin
        _T_136_15 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h10 == auto_in_a_bits_source) begin
        _T_136_16 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h11 == auto_in_a_bits_source) begin
        _T_136_17 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h12 == auto_in_a_bits_source) begin
        _T_136_18 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h13 == auto_in_a_bits_source) begin
        _T_136_19 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h14 == auto_in_a_bits_source) begin
        _T_136_20 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h15 == auto_in_a_bits_source) begin
        _T_136_21 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h16 == auto_in_a_bits_source) begin
        _T_136_22 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h17 == auto_in_a_bits_source) begin
        _T_136_23 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h18 == auto_in_a_bits_source) begin
        _T_136_24 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h19 == auto_in_a_bits_source) begin
        _T_136_25 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h1a == auto_in_a_bits_source) begin
        _T_136_26 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h1b == auto_in_a_bits_source) begin
        _T_136_27 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h1c == auto_in_a_bits_source) begin
        _T_136_28 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h1d == auto_in_a_bits_source) begin
        _T_136_29 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h1e == auto_in_a_bits_source) begin
        _T_136_30 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h1f == auto_in_a_bits_source) begin
        _T_136_31 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h20 == auto_in_a_bits_source) begin
        _T_136_32 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h21 == auto_in_a_bits_source) begin
        _T_136_33 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h22 == auto_in_a_bits_source) begin
        _T_136_34 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h23 == auto_in_a_bits_source) begin
        _T_136_35 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h24 == auto_in_a_bits_source) begin
        _T_136_36 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h25 == auto_in_a_bits_source) begin
        _T_136_37 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h26 == auto_in_a_bits_source) begin
        _T_136_38 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h27 == auto_in_a_bits_source) begin
        _T_136_39 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h28 == auto_in_a_bits_source) begin
        _T_136_40 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h29 == auto_in_a_bits_source) begin
        _T_136_41 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h2a == auto_in_a_bits_source) begin
        _T_136_42 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h2b == auto_in_a_bits_source) begin
        _T_136_43 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h2c == auto_in_a_bits_source) begin
        _T_136_44 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h2d == auto_in_a_bits_source) begin
        _T_136_45 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h2e == auto_in_a_bits_source) begin
        _T_136_46 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h2f == auto_in_a_bits_source) begin
        _T_136_47 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h30 == auto_in_a_bits_source) begin
        _T_136_48 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h31 == auto_in_a_bits_source) begin
        _T_136_49 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h32 == auto_in_a_bits_source) begin
        _T_136_50 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h33 == auto_in_a_bits_source) begin
        _T_136_51 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h34 == auto_in_a_bits_source) begin
        _T_136_52 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h35 == auto_in_a_bits_source) begin
        _T_136_53 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h36 == auto_in_a_bits_source) begin
        _T_136_54 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h37 == auto_in_a_bits_source) begin
        _T_136_55 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h38 == auto_in_a_bits_source) begin
        _T_136_56 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h39 == auto_in_a_bits_source) begin
        _T_136_57 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h3a == auto_in_a_bits_source) begin
        _T_136_58 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h3b == auto_in_a_bits_source) begin
        _T_136_59 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h3c == auto_in_a_bits_source) begin
        _T_136_60 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h3d == auto_in_a_bits_source) begin
        _T_136_61 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h3e == auto_in_a_bits_source) begin
        _T_136_62 <= _T_50;
      end
    end
    if (_T_30) begin
      if (6'h3f == auto_in_a_bits_source) begin
        _T_136_63 <= _T_50;
      end
    end
    if (_T_129) begin
      if (6'h3f == _T_118_bits_source) begin
        _T_141 <= _T_136_63;
      end else begin
        if (6'h3e == _T_118_bits_source) begin
          _T_141 <= _T_136_62;
        end else begin
          if (6'h3d == _T_118_bits_source) begin
            _T_141 <= _T_136_61;
          end else begin
            if (6'h3c == _T_118_bits_source) begin
              _T_141 <= _T_136_60;
            end else begin
              if (6'h3b == _T_118_bits_source) begin
                _T_141 <= _T_136_59;
              end else begin
                if (6'h3a == _T_118_bits_source) begin
                  _T_141 <= _T_136_58;
                end else begin
                  if (6'h39 == _T_118_bits_source) begin
                    _T_141 <= _T_136_57;
                  end else begin
                    if (6'h38 == _T_118_bits_source) begin
                      _T_141 <= _T_136_56;
                    end else begin
                      if (6'h37 == _T_118_bits_source) begin
                        _T_141 <= _T_136_55;
                      end else begin
                        if (6'h36 == _T_118_bits_source) begin
                          _T_141 <= _T_136_54;
                        end else begin
                          if (6'h35 == _T_118_bits_source) begin
                            _T_141 <= _T_136_53;
                          end else begin
                            if (6'h34 == _T_118_bits_source) begin
                              _T_141 <= _T_136_52;
                            end else begin
                              if (6'h33 == _T_118_bits_source) begin
                                _T_141 <= _T_136_51;
                              end else begin
                                if (6'h32 == _T_118_bits_source) begin
                                  _T_141 <= _T_136_50;
                                end else begin
                                  if (6'h31 == _T_118_bits_source) begin
                                    _T_141 <= _T_136_49;
                                  end else begin
                                    if (6'h30 == _T_118_bits_source) begin
                                      _T_141 <= _T_136_48;
                                    end else begin
                                      if (6'h2f == _T_118_bits_source) begin
                                        _T_141 <= _T_136_47;
                                      end else begin
                                        if (6'h2e == _T_118_bits_source) begin
                                          _T_141 <= _T_136_46;
                                        end else begin
                                          if (6'h2d == _T_118_bits_source) begin
                                            _T_141 <= _T_136_45;
                                          end else begin
                                            if (6'h2c == _T_118_bits_source) begin
                                              _T_141 <= _T_136_44;
                                            end else begin
                                              if (6'h2b == _T_118_bits_source) begin
                                                _T_141 <= _T_136_43;
                                              end else begin
                                                if (6'h2a == _T_118_bits_source) begin
                                                  _T_141 <= _T_136_42;
                                                end else begin
                                                  if (6'h29 == _T_118_bits_source) begin
                                                    _T_141 <= _T_136_41;
                                                  end else begin
                                                    if (6'h28 == _T_118_bits_source) begin
                                                      _T_141 <= _T_136_40;
                                                    end else begin
                                                      if (6'h27 == _T_118_bits_source) begin
                                                        _T_141 <= _T_136_39;
                                                      end else begin
                                                        if (6'h26 == _T_118_bits_source) begin
                                                          _T_141 <= _T_136_38;
                                                        end else begin
                                                          if (6'h25 == _T_118_bits_source) begin
                                                            _T_141 <= _T_136_37;
                                                          end else begin
                                                            if (6'h24 == _T_118_bits_source) begin
                                                              _T_141 <= _T_136_36;
                                                            end else begin
                                                              if (6'h23 == _T_118_bits_source) begin
                                                                _T_141 <= _T_136_35;
                                                              end else begin
                                                                if (6'h22 == _T_118_bits_source) begin
                                                                  _T_141 <= _T_136_34;
                                                                end else begin
                                                                  if (6'h21 == _T_118_bits_source) begin
                                                                    _T_141 <= _T_136_33;
                                                                  end else begin
                                                                    if (6'h20 == _T_118_bits_source) begin
                                                                      _T_141 <= _T_136_32;
                                                                    end else begin
                                                                      if (6'h1f == _T_118_bits_source) begin
                                                                        _T_141 <= _T_136_31;
                                                                      end else begin
                                                                        if (6'h1e == _T_118_bits_source) begin
                                                                          _T_141 <= _T_136_30;
                                                                        end else begin
                                                                          if (6'h1d == _T_118_bits_source) begin
                                                                            _T_141 <= _T_136_29;
                                                                          end else begin
                                                                            if (6'h1c == _T_118_bits_source) begin
                                                                              _T_141 <= _T_136_28;
                                                                            end else begin
                                                                              if (6'h1b == _T_118_bits_source) begin
                                                                                _T_141 <= _T_136_27;
                                                                              end else begin
                                                                                if (6'h1a == _T_118_bits_source) begin
                                                                                  _T_141 <= _T_136_26;
                                                                                end else begin
                                                                                  if (6'h19 == _T_118_bits_source) begin
                                                                                    _T_141 <= _T_136_25;
                                                                                  end else begin
                                                                                    if (6'h18 == _T_118_bits_source) begin
                                                                                      _T_141 <= _T_136_24;
                                                                                    end else begin
                                                                                      if (6'h17 == _T_118_bits_source) begin
                                                                                        _T_141 <= _T_136_23;
                                                                                      end else begin
                                                                                        if (6'h16 == _T_118_bits_source) begin
                                                                                          _T_141 <= _T_136_22;
                                                                                        end else begin
                                                                                          if (6'h15 == _T_118_bits_source) begin
                                                                                            _T_141 <= _T_136_21;
                                                                                          end else begin
                                                                                            if (6'h14 == _T_118_bits_source) begin
                                                                                              _T_141 <= _T_136_20;
                                                                                            end else begin
                                                                                              if (6'h13 == _T_118_bits_source) begin
                                                                                                _T_141 <= _T_136_19;
                                                                                              end else begin
                                                                                                if (6'h12 == _T_118_bits_source) begin
                                                                                                  _T_141 <= _T_136_18;
                                                                                                end else begin
                                                                                                  if (6'h11 == _T_118_bits_source) begin
                                                                                                    _T_141 <= _T_136_17;
                                                                                                  end else begin
                                                                                                    if (6'h10 == _T_118_bits_source) begin
                                                                                                      _T_141 <= _T_136_16;
                                                                                                    end else begin
                                                                                                      if (6'hf == _T_118_bits_source) begin
                                                                                                        _T_141 <= _T_136_15;
                                                                                                      end else begin
                                                                                                        if (6'he == _T_118_bits_source) begin
                                                                                                          _T_141 <= _T_136_14;
                                                                                                        end else begin
                                                                                                          if (6'hd == _T_118_bits_source) begin
                                                                                                            _T_141 <= _T_136_13;
                                                                                                          end else begin
                                                                                                            if (6'hc == _T_118_bits_source) begin
                                                                                                              _T_141 <= _T_136_12;
                                                                                                            end else begin
                                                                                                              if (6'hb == _T_118_bits_source) begin
                                                                                                                _T_141 <= _T_136_11;
                                                                                                              end else begin
                                                                                                                if (6'ha == _T_118_bits_source) begin
                                                                                                                  _T_141 <= _T_136_10;
                                                                                                                end else begin
                                                                                                                  if (6'h9 == _T_118_bits_source) begin
                                                                                                                    _T_141 <= _T_136_9;
                                                                                                                  end else begin
                                                                                                                    if (6'h8 == _T_118_bits_source) begin
                                                                                                                      _T_141 <= _T_136_8;
                                                                                                                    end else begin
                                                                                                                      if (6'h7 == _T_118_bits_source) begin
                                                                                                                        _T_141 <= _T_136_7;
                                                                                                                      end else begin
                                                                                                                        if (6'h6 == _T_118_bits_source) begin
                                                                                                                          _T_141 <= _T_136_6;
                                                                                                                        end else begin
                                                                                                                          if (6'h5 == _T_118_bits_source) begin
                                                                                                                            _T_141 <= _T_136_5;
                                                                                                                          end else begin
                                                                                                                            if (6'h4 == _T_118_bits_source) begin
                                                                                                                              _T_141 <= _T_136_4;
                                                                                                                            end else begin
                                                                                                                              if (6'h3 == _T_118_bits_source) begin
                                                                                                                                _T_141 <= _T_136_3;
                                                                                                                              end else begin
                                                                                                                                if (6'h2 == _T_118_bits_source) begin
                                                                                                                                  _T_141 <= _T_136_2;
                                                                                                                                end else begin
                                                                                                                                  if (6'h1 == _T_118_bits_source) begin
                                                                                                                                    _T_141 <= _T_136_1;
                                                                                                                                  end else begin
                                                                                                                                    _T_141 <= _T_136_0;
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_182 <= 1'h0;
    end else begin
      if (_T_197) begin
        if (_T_186) begin
          _T_182 <= 1'h0;
        end else begin
          _T_182 <= _T_199;
        end
      end
    end
    if (reset) begin
      _T_195 <= 1'h0;
    end else begin
      if (_T_197) begin
        if (_T_186) begin
          _T_195 <= 1'h0;
        end else begin
          _T_195 <= _T_196;
        end
      end
    end
  end
endmodule
module dual_TLWidthWidget_2( 
  input         clock, 
  input         reset, 
  output        auto_in_a_ready, 
  input         auto_in_a_valid, 
  input  [2:0]  auto_in_a_bits_opcode, 
  input  [2:0]  auto_in_a_bits_param, 
  input  [2:0]  auto_in_a_bits_size, 
  input  [6:0]  auto_in_a_bits_source, 
  input  [28:0] auto_in_a_bits_address, 
  input  [7:0]  auto_in_a_bits_mask, 
  input         auto_in_a_bits_corrupt, 
  output        auto_in_c_ready, 
  input         auto_in_c_valid, 
  input  [2:0]  auto_in_c_bits_opcode, 
  input  [2:0]  auto_in_c_bits_param, 
  input  [2:0]  auto_in_c_bits_size, 
  input  [6:0]  auto_in_c_bits_source, 
  input  [28:0] auto_in_c_bits_address, 
  input         auto_in_c_bits_corrupt, 
  input         auto_in_d_ready, 
  output        auto_in_d_valid, 
  output [2:0]  auto_in_d_bits_opcode, 
  output [1:0]  auto_in_d_bits_param, 
  output [2:0]  auto_in_d_bits_size, 
  output [6:0]  auto_in_d_bits_source, 
  output        auto_in_d_bits_sink, 
  output        auto_in_d_bits_denied, 
  output [63:0] auto_in_d_bits_data, 
  output        auto_in_d_bits_corrupt, 
  input         auto_in_e_valid, 
  input         auto_out_a_ready, 
  output        auto_out_a_valid, 
  output [2:0]  auto_out_a_bits_opcode, 
  output [2:0]  auto_out_a_bits_param, 
  output [2:0]  auto_out_a_bits_size, 
  output [6:0]  auto_out_a_bits_source, 
  output [28:0] auto_out_a_bits_address, 
  output [3:0]  auto_out_a_bits_mask, 
  output        auto_out_a_bits_corrupt, 
  input         auto_out_c_ready, 
  output        auto_out_c_valid, 
  output [2:0]  auto_out_c_bits_opcode, 
  output [2:0]  auto_out_c_bits_param, 
  output [2:0]  auto_out_c_bits_size, 
  output [6:0]  auto_out_c_bits_source, 
  output [28:0] auto_out_c_bits_address, 
  output        auto_out_c_bits_corrupt, 
  output        auto_out_d_ready, 
  input         auto_out_d_valid, 
  input  [2:0]  auto_out_d_bits_opcode, 
  input  [1:0]  auto_out_d_bits_param, 
  input  [2:0]  auto_out_d_bits_size, 
  input  [6:0]  auto_out_d_bits_source, 
  input         auto_out_d_bits_sink, 
  input         auto_out_d_bits_denied, 
  input  [31:0] auto_out_d_bits_data, 
  input         auto_out_d_bits_corrupt, 
  output        auto_out_e_valid 
);
  wire  TLMonitor_clock; 
  wire  TLMonitor_reset; 
  wire  TLMonitor_io_in_a_ready; 
  wire  TLMonitor_io_in_a_valid; 
  wire [2:0] TLMonitor_io_in_a_bits_opcode; 
  wire [2:0] TLMonitor_io_in_a_bits_param; 
  wire [2:0] TLMonitor_io_in_a_bits_size; 
  wire [6:0] TLMonitor_io_in_a_bits_source; 
  wire [28:0] TLMonitor_io_in_a_bits_address; 
  wire [7:0] TLMonitor_io_in_a_bits_mask; 
  wire  TLMonitor_io_in_a_bits_corrupt; 
  wire  TLMonitor_io_in_c_ready; 
  wire  TLMonitor_io_in_c_valid; 
  wire [2:0] TLMonitor_io_in_c_bits_opcode; 
  wire [2:0] TLMonitor_io_in_c_bits_param; 
  wire [2:0] TLMonitor_io_in_c_bits_size; 
  wire [6:0] TLMonitor_io_in_c_bits_source; 
  wire [28:0] TLMonitor_io_in_c_bits_address; 
  wire  TLMonitor_io_in_c_bits_corrupt; 
  wire  TLMonitor_io_in_d_ready; 
  wire  TLMonitor_io_in_d_valid; 
  wire [2:0] TLMonitor_io_in_d_bits_opcode; 
  wire [1:0] TLMonitor_io_in_d_bits_param; 
  wire [2:0] TLMonitor_io_in_d_bits_size; 
  wire [6:0] TLMonitor_io_in_d_bits_source; 
  wire  TLMonitor_io_in_d_bits_sink; 
  wire  TLMonitor_io_in_d_bits_denied; 
  wire  TLMonitor_io_in_d_bits_corrupt; 
  wire  TLMonitor_io_in_e_valid; 
  wire  Repeater_clock; 
  wire  Repeater_reset; 
  wire  Repeater_io_repeat; 
  wire  Repeater_io_enq_ready; 
  wire  Repeater_io_enq_valid; 
  wire [2:0] Repeater_io_enq_bits_opcode; 
  wire [2:0] Repeater_io_enq_bits_param; 
  wire [2:0] Repeater_io_enq_bits_size; 
  wire [6:0] Repeater_io_enq_bits_source; 
  wire [28:0] Repeater_io_enq_bits_address; 
  wire [7:0] Repeater_io_enq_bits_mask; 
  wire  Repeater_io_enq_bits_corrupt; 
  wire  Repeater_io_deq_ready; 
  wire  Repeater_io_deq_valid; 
  wire [2:0] Repeater_io_deq_bits_opcode; 
  wire [2:0] Repeater_io_deq_bits_param; 
  wire [2:0] Repeater_io_deq_bits_size; 
  wire [6:0] Repeater_io_deq_bits_source; 
  wire [28:0] Repeater_io_deq_bits_address; 
  wire [7:0] Repeater_io_deq_bits_mask; 
  wire  Repeater_io_deq_bits_corrupt; 
  wire  Repeater_1_clock; 
  wire  Repeater_1_reset; 
  wire  Repeater_1_io_repeat; 
  wire  Repeater_1_io_enq_ready; 
  wire  Repeater_1_io_enq_valid; 
  wire [2:0] Repeater_1_io_enq_bits_opcode; 
  wire [2:0] Repeater_1_io_enq_bits_param; 
  wire [2:0] Repeater_1_io_enq_bits_size; 
  wire [6:0] Repeater_1_io_enq_bits_source; 
  wire [28:0] Repeater_1_io_enq_bits_address; 
  wire  Repeater_1_io_enq_bits_corrupt; 
  wire  Repeater_1_io_deq_ready; 
  wire  Repeater_1_io_deq_valid; 
  wire [2:0] Repeater_1_io_deq_bits_opcode; 
  wire [2:0] Repeater_1_io_deq_bits_param; 
  wire [2:0] Repeater_1_io_deq_bits_size; 
  wire [6:0] Repeater_1_io_deq_bits_source; 
  wire [28:0] Repeater_1_io_deq_bits_address; 
  wire  Repeater_1_io_deq_bits_corrupt; 
  wire [2:0] _T_9_bits_opcode; 
  wire  _T_13; 
  wire  _T_14; 
  wire [2:0] _T_9_bits_size; 
  wire [9:0] _T_16; 
  wire [2:0] _T_17; 
  wire [2:0] _T_18; 
  wire  _T_19; 
  reg  _T_20; 
  reg [31:0] _RAND_0;
  wire  _T_22; 
  wire  _T_23; 
  wire  _T_24; 
  wire  _T_9_valid; 
  wire  _T_25; 
  wire  _T_27; 
  wire [28:0] _T_9_bits_address; 
  wire  _T_28; 
  wire  _T_29; 
  wire [7:0] _T_9_bits_mask; 
  wire [3:0] _T_33; 
  wire [3:0] _T_34; 
  wire  _T_37; 
  wire [9:0] _T_39; 
  wire [2:0] _T_40; 
  wire [2:0] _T_41; 
  wire  _T_42; 
  reg  _T_43; 
  reg [31:0] _RAND_1;
  wire  _T_45; 
  wire  _T_46; 
  wire  _T_47; 
  wire  _T_49; 
  wire  _T_51; 
  reg  _T_56; 
  reg [31:0] _RAND_2;
  wire  _T_57; 
  wire  _T_61; 
  wire  _T_62; 
  wire  _T_58; 
  wire  _T_60; 
  reg [31:0] _T_64_0; 
  reg [31:0] _RAND_3;
  wire [31:0] _T_65; 
  wire  _T_69; 
  wire [2:0] _T_174_bits_opcode; 
  wire  _T_178; 
  wire [2:0] _T_174_bits_size; 
  wire [9:0] _T_180; 
  wire [2:0] _T_181; 
  wire [2:0] _T_182; 
  wire  _T_183; 
  reg  _T_184; 
  reg [31:0] _RAND_4;
  wire  _T_186; 
  wire  _T_187; 
  wire  _T_188; 
  wire  _T_174_valid; 
  wire  _T_189; 
  wire  _T_191; 
  dual_TLMonitor_18 dual_TLMonitor ( 
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_io_in_a_bits_corrupt),
    .io_in_c_ready(TLMonitor_io_in_c_ready),
    .io_in_c_valid(TLMonitor_io_in_c_valid),
    .io_in_c_bits_opcode(TLMonitor_io_in_c_bits_opcode),
    .io_in_c_bits_param(TLMonitor_io_in_c_bits_param),
    .io_in_c_bits_size(TLMonitor_io_in_c_bits_size),
    .io_in_c_bits_source(TLMonitor_io_in_c_bits_source),
    .io_in_c_bits_address(TLMonitor_io_in_c_bits_address),
    .io_in_c_bits_corrupt(TLMonitor_io_in_c_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt),
    .io_in_e_valid(TLMonitor_io_in_e_valid)
  );
  dual_Repeater_4 dual_Repeater_top ( 
    .clock(Repeater_clock),
    .reset(Repeater_reset),
    .io_repeat(Repeater_io_repeat),
    .io_enq_ready(Repeater_io_enq_ready),
    .io_enq_valid(Repeater_io_enq_valid),
    .io_enq_bits_opcode(Repeater_io_enq_bits_opcode),
    .io_enq_bits_param(Repeater_io_enq_bits_param),
    .io_enq_bits_size(Repeater_io_enq_bits_size),
    .io_enq_bits_source(Repeater_io_enq_bits_source),
    .io_enq_bits_address(Repeater_io_enq_bits_address),
    .io_enq_bits_mask(Repeater_io_enq_bits_mask),
    .io_enq_bits_corrupt(Repeater_io_enq_bits_corrupt),
    .io_deq_ready(Repeater_io_deq_ready),
    .io_deq_valid(Repeater_io_deq_valid),
    .io_deq_bits_opcode(Repeater_io_deq_bits_opcode),
    .io_deq_bits_param(Repeater_io_deq_bits_param),
    .io_deq_bits_size(Repeater_io_deq_bits_size),
    .io_deq_bits_source(Repeater_io_deq_bits_source),
    .io_deq_bits_address(Repeater_io_deq_bits_address),
    .io_deq_bits_mask(Repeater_io_deq_bits_mask),
    .io_deq_bits_corrupt(Repeater_io_deq_bits_corrupt)
  );
  dual_Repeater_5 dual_Repeater_1 ( 
    .clock(Repeater_1_clock),
    .reset(Repeater_1_reset),
    .io_repeat(Repeater_1_io_repeat),
    .io_enq_ready(Repeater_1_io_enq_ready),
    .io_enq_valid(Repeater_1_io_enq_valid),
    .io_enq_bits_opcode(Repeater_1_io_enq_bits_opcode),
    .io_enq_bits_param(Repeater_1_io_enq_bits_param),
    .io_enq_bits_size(Repeater_1_io_enq_bits_size),
    .io_enq_bits_source(Repeater_1_io_enq_bits_source),
    .io_enq_bits_address(Repeater_1_io_enq_bits_address),
    .io_enq_bits_corrupt(Repeater_1_io_enq_bits_corrupt),
    .io_deq_ready(Repeater_1_io_deq_ready),
    .io_deq_valid(Repeater_1_io_deq_valid),
    .io_deq_bits_opcode(Repeater_1_io_deq_bits_opcode),
    .io_deq_bits_param(Repeater_1_io_deq_bits_param),
    .io_deq_bits_size(Repeater_1_io_deq_bits_size),
    .io_deq_bits_source(Repeater_1_io_deq_bits_source),
    .io_deq_bits_address(Repeater_1_io_deq_bits_address),
    .io_deq_bits_corrupt(Repeater_1_io_deq_bits_corrupt)
  );
  assign _T_9_bits_opcode = Repeater_io_deq_bits_opcode; 
  assign _T_13 = _T_9_bits_opcode[2]; 
  assign _T_14 = _T_13 == 1'h0; 
  assign _T_9_bits_size = Repeater_io_deq_bits_size; 
  assign _T_16 = 10'h7 << _T_9_bits_size; 
  assign _T_17 = _T_16[2:0]; 
  assign _T_18 = ~ _T_17; 
  assign _T_19 = _T_18[2:2]; 
  assign _T_22 = _T_20 == _T_19; 
  assign _T_23 = _T_14 == 1'h0; 
  assign _T_24 = _T_22 | _T_23; 
  assign _T_9_valid = Repeater_io_deq_valid; 
  assign _T_25 = auto_out_a_ready & _T_9_valid; 
  assign _T_27 = _T_20 + 1'h1; 
  assign _T_9_bits_address = Repeater_io_deq_bits_address; 
  assign _T_28 = _T_9_bits_address[2]; 
  assign _T_29 = _T_28 | _T_20; 
  assign _T_9_bits_mask = Repeater_io_deq_bits_mask; 
  assign _T_33 = _T_9_bits_mask[3:0]; 
  assign _T_34 = _T_9_bits_mask[7:4]; 
  assign _T_37 = auto_out_d_bits_opcode[0]; 
  assign _T_39 = 10'h7 << auto_out_d_bits_size; 
  assign _T_40 = _T_39[2:0]; 
  assign _T_41 = ~ _T_40; 
  assign _T_42 = _T_41[2:2]; 
  assign _T_45 = _T_43 == _T_42; 
  assign _T_46 = _T_37 == 1'h0; 
  assign _T_47 = _T_45 | _T_46; 
  assign _T_49 = _T_43 & _T_42; 
  assign _T_51 = _T_49 == 1'h0; 
  assign _T_57 = auto_out_d_bits_corrupt | _T_56; 
  assign _T_61 = _T_47 == 1'h0; 
  assign _T_62 = auto_in_d_ready | _T_61; 
  assign _T_58 = _T_62 & auto_out_d_valid; 
  assign _T_60 = _T_43 + 1'h1; 
  assign _T_65 = _T_51 ? auto_out_d_bits_data : _T_64_0; 
  assign _T_69 = _T_58 & _T_61; 
  assign _T_174_bits_opcode = Repeater_1_io_deq_bits_opcode; 
  assign _T_178 = _T_174_bits_opcode[0]; 
  assign _T_174_bits_size = Repeater_1_io_deq_bits_size; 
  assign _T_180 = 10'h7 << _T_174_bits_size; 
  assign _T_181 = _T_180[2:0]; 
  assign _T_182 = ~ _T_181; 
  assign _T_183 = _T_182[2:2]; 
  assign _T_186 = _T_184 == _T_183; 
  assign _T_187 = _T_178 == 1'h0; 
  assign _T_188 = _T_186 | _T_187; 
  assign _T_174_valid = Repeater_1_io_deq_valid; 
  assign _T_189 = auto_out_c_ready & _T_174_valid; 
  assign _T_191 = _T_184 + 1'h1; 
  assign auto_in_a_ready = Repeater_io_enq_ready; 
  assign auto_in_c_ready = Repeater_1_io_enq_ready; 
  assign auto_in_d_valid = auto_out_d_valid & _T_47; 
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; 
  assign auto_in_d_bits_param = auto_out_d_bits_param; 
  assign auto_in_d_bits_size = auto_out_d_bits_size; 
  assign auto_in_d_bits_source = auto_out_d_bits_source; 
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; 
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; 
  assign auto_in_d_bits_data = {auto_out_d_bits_data,_T_65}; 
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt | _T_56; 
  assign auto_out_a_valid = Repeater_io_deq_valid; 
  assign auto_out_a_bits_opcode = Repeater_io_deq_bits_opcode; 
  assign auto_out_a_bits_param = Repeater_io_deq_bits_param; 
  assign auto_out_a_bits_size = Repeater_io_deq_bits_size; 
  assign auto_out_a_bits_source = Repeater_io_deq_bits_source; 
  assign auto_out_a_bits_address = Repeater_io_deq_bits_address; 
  assign auto_out_a_bits_mask = _T_29 ? _T_34 : _T_33; 
  assign auto_out_a_bits_corrupt = Repeater_io_deq_bits_corrupt; 
  assign auto_out_c_valid = Repeater_1_io_deq_valid; 
  assign auto_out_c_bits_opcode = Repeater_1_io_deq_bits_opcode; 
  assign auto_out_c_bits_param = Repeater_1_io_deq_bits_param; 
  assign auto_out_c_bits_size = Repeater_1_io_deq_bits_size; 
  assign auto_out_c_bits_source = Repeater_1_io_deq_bits_source; 
  assign auto_out_c_bits_address = Repeater_1_io_deq_bits_address; 
  assign auto_out_c_bits_corrupt = Repeater_1_io_deq_bits_corrupt; 
  assign auto_out_d_ready = auto_in_d_ready | _T_61; 
  assign auto_out_e_valid = auto_in_e_valid; 
  assign TLMonitor_clock = clock; 
  assign TLMonitor_reset = reset; 
  assign TLMonitor_io_in_a_ready = Repeater_io_enq_ready; 
  assign TLMonitor_io_in_a_valid = auto_in_a_valid; 
  assign TLMonitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; 
  assign TLMonitor_io_in_a_bits_param = auto_in_a_bits_param; 
  assign TLMonitor_io_in_a_bits_size = auto_in_a_bits_size; 
  assign TLMonitor_io_in_a_bits_source = auto_in_a_bits_source; 
  assign TLMonitor_io_in_a_bits_address = auto_in_a_bits_address; 
  assign TLMonitor_io_in_a_bits_mask = auto_in_a_bits_mask; 
  assign TLMonitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; 
  assign TLMonitor_io_in_c_ready = Repeater_1_io_enq_ready; 
  assign TLMonitor_io_in_c_valid = auto_in_c_valid; 
  assign TLMonitor_io_in_c_bits_opcode = auto_in_c_bits_opcode; 
  assign TLMonitor_io_in_c_bits_param = auto_in_c_bits_param; 
  assign TLMonitor_io_in_c_bits_size = auto_in_c_bits_size; 
  assign TLMonitor_io_in_c_bits_source = auto_in_c_bits_source; 
  assign TLMonitor_io_in_c_bits_address = auto_in_c_bits_address; 
  assign TLMonitor_io_in_c_bits_corrupt = auto_in_c_bits_corrupt; 
  assign TLMonitor_io_in_d_ready = auto_in_d_ready; 
  assign TLMonitor_io_in_d_valid = auto_out_d_valid & _T_47; 
  assign TLMonitor_io_in_d_bits_opcode = auto_out_d_bits_opcode; 
  assign TLMonitor_io_in_d_bits_param = auto_out_d_bits_param; 
  assign TLMonitor_io_in_d_bits_size = auto_out_d_bits_size; 
  assign TLMonitor_io_in_d_bits_source = auto_out_d_bits_source; 
  assign TLMonitor_io_in_d_bits_sink = auto_out_d_bits_sink; 
  assign TLMonitor_io_in_d_bits_denied = auto_out_d_bits_denied; 
  assign TLMonitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt | _T_56; 
  assign TLMonitor_io_in_e_valid = auto_in_e_valid; 
  assign Repeater_clock = clock; 
  assign Repeater_reset = reset; 
  assign Repeater_io_repeat = _T_24 == 1'h0; 
  assign Repeater_io_enq_valid = auto_in_a_valid; 
  assign Repeater_io_enq_bits_opcode = auto_in_a_bits_opcode; 
  assign Repeater_io_enq_bits_param = auto_in_a_bits_param; 
  assign Repeater_io_enq_bits_size = auto_in_a_bits_size; 
  assign Repeater_io_enq_bits_source = auto_in_a_bits_source; 
  assign Repeater_io_enq_bits_address = auto_in_a_bits_address; 
  assign Repeater_io_enq_bits_mask = auto_in_a_bits_mask; 
  assign Repeater_io_enq_bits_corrupt = auto_in_a_bits_corrupt; 
  assign Repeater_io_deq_ready = auto_out_a_ready; 
  assign Repeater_1_clock = clock; 
  assign Repeater_1_reset = reset; 
  assign Repeater_1_io_repeat = _T_188 == 1'h0; 
  assign Repeater_1_io_enq_valid = auto_in_c_valid; 
  assign Repeater_1_io_enq_bits_opcode = auto_in_c_bits_opcode; 
  assign Repeater_1_io_enq_bits_param = auto_in_c_bits_param; 
  assign Repeater_1_io_enq_bits_size = auto_in_c_bits_size; 
  assign Repeater_1_io_enq_bits_source = auto_in_c_bits_source; 
  assign Repeater_1_io_enq_bits_address = auto_in_c_bits_address; 
  assign Repeater_1_io_enq_bits_corrupt = auto_in_c_bits_corrupt; 
  assign Repeater_1_io_deq_ready = auto_out_c_ready; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_20 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_43 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_56 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_64_0 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_184 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_20 <= 1'h0;
    end else begin
      if (_T_25) begin
        if (_T_24) begin
          _T_20 <= 1'h0;
        end else begin
          _T_20 <= _T_27;
        end
      end
    end
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      if (_T_58) begin
        if (_T_47) begin
          _T_43 <= 1'h0;
        end else begin
          _T_43 <= _T_60;
        end
      end
    end
    if (reset) begin
      _T_56 <= 1'h0;
    end else begin
      if (_T_58) begin
        if (_T_47) begin
          _T_56 <= 1'h0;
        end else begin
          _T_56 <= _T_57;
        end
      end
    end
    if (_T_69) begin
      if (_T_51) begin
        _T_64_0 <= auto_out_d_bits_data;
      end
    end
    if (reset) begin
      _T_184 <= 1'h0;
    end else begin
      if (_T_189) begin
        if (_T_188) begin
          _T_184 <= 1'h0;
        end else begin
          _T_184 <= _T_191;
        end
      end
    end
  end
endmodule
module dual_TLWidthWidget( 
  input         clock, 
  input         reset, 
  output        auto_in_a_ready, 
  input         auto_in_a_valid, 
  input  [2:0]  auto_in_a_bits_opcode, 
  input  [2:0]  auto_in_a_bits_param, 
  input  [2:0]  auto_in_a_bits_size, 
  input  [2:0]  auto_in_a_bits_source, 
  input  [31:0] auto_in_a_bits_address, 
  input  [7:0]  auto_in_a_bits_mask, 
  input  [63:0] auto_in_a_bits_data, 
  input         auto_in_a_bits_corrupt, 
  input         auto_in_d_ready, 
  output        auto_in_d_valid, 
  output [2:0]  auto_in_d_bits_opcode, 
  output [2:0]  auto_in_d_bits_size, 
  output [2:0]  auto_in_d_bits_source, 
  output        auto_in_d_bits_denied, 
  output [63:0] auto_in_d_bits_data, 
  output        auto_in_d_bits_corrupt, 
  input         auto_out_a_ready, 
  output        auto_out_a_valid, 
  output [2:0]  auto_out_a_bits_opcode, 
  output [2:0]  auto_out_a_bits_param, 
  output [2:0]  auto_out_a_bits_size, 
  output [2:0]  auto_out_a_bits_source, 
  output [31:0] auto_out_a_bits_address, 
  output [3:0]  auto_out_a_bits_mask, 
  output [31:0] auto_out_a_bits_data, 
  output        auto_out_a_bits_corrupt, 
  output        auto_out_d_ready, 
  input         auto_out_d_valid, 
  input  [2:0]  auto_out_d_bits_opcode, 
  input  [1:0]  auto_out_d_bits_param, 
  input  [2:0]  auto_out_d_bits_size, 
  input  [2:0]  auto_out_d_bits_source, 
  input  [5:0]  auto_out_d_bits_sink, 
  input         auto_out_d_bits_denied, 
  input  [31:0] auto_out_d_bits_data, 
  input         auto_out_d_bits_corrupt 
);
  wire  TLMonitor_clock; 
  wire  TLMonitor_reset; 
  wire  TLMonitor_io_in_a_ready; 
  wire  TLMonitor_io_in_a_valid; 
  wire [2:0] TLMonitor_io_in_a_bits_opcode; 
  wire [2:0] TLMonitor_io_in_a_bits_param; 
  wire [2:0] TLMonitor_io_in_a_bits_size; 
  wire [2:0] TLMonitor_io_in_a_bits_source; 
  wire [31:0] TLMonitor_io_in_a_bits_address; 
  wire [7:0] TLMonitor_io_in_a_bits_mask; 
  wire  TLMonitor_io_in_a_bits_corrupt; 
  wire  TLMonitor_io_in_d_ready; 
  wire  TLMonitor_io_in_d_valid; 
  wire [2:0] TLMonitor_io_in_d_bits_opcode; 
  wire [1:0] TLMonitor_io_in_d_bits_param; 
  wire [2:0] TLMonitor_io_in_d_bits_size; 
  wire [2:0] TLMonitor_io_in_d_bits_source; 
  wire [5:0] TLMonitor_io_in_d_bits_sink; 
  wire  TLMonitor_io_in_d_bits_denied; 
  wire  TLMonitor_io_in_d_bits_corrupt; 
  wire  Repeater_clock; 
  wire  Repeater_reset; 
  wire  Repeater_io_repeat; 
  wire  Repeater_io_enq_ready; 
  wire  Repeater_io_enq_valid; 
  wire [2:0] Repeater_io_enq_bits_opcode; 
  wire [2:0] Repeater_io_enq_bits_param; 
  wire [2:0] Repeater_io_enq_bits_size; 
  wire [2:0] Repeater_io_enq_bits_source; 
  wire [31:0] Repeater_io_enq_bits_address; 
  wire [7:0] Repeater_io_enq_bits_mask; 
  wire [63:0] Repeater_io_enq_bits_data; 
  wire  Repeater_io_enq_bits_corrupt; 
  wire  Repeater_io_deq_ready; 
  wire  Repeater_io_deq_valid; 
  wire [2:0] Repeater_io_deq_bits_opcode; 
  wire [2:0] Repeater_io_deq_bits_param; 
  wire [2:0] Repeater_io_deq_bits_size; 
  wire [2:0] Repeater_io_deq_bits_source; 
  wire [31:0] Repeater_io_deq_bits_address; 
  wire [7:0] Repeater_io_deq_bits_mask; 
  wire [63:0] Repeater_io_deq_bits_data; 
  wire  Repeater_io_deq_bits_corrupt; 
  wire [31:0] _T_10; 
  wire [31:0] _T_11; 
  wire [63:0] _T_12; 
  wire [2:0] _T_9_bits_opcode; 
  wire  _T_13; 
  wire  _T_14; 
  wire [2:0] _T_9_bits_size; 
  wire [9:0] _T_16; 
  wire [2:0] _T_17; 
  wire [2:0] _T_18; 
  wire  _T_19; 
  reg  _T_20; 
  reg [31:0] _RAND_0;
  wire  _T_22; 
  wire  _T_23; 
  wire  _T_24; 
  wire  _T_9_valid; 
  wire  _T_25; 
  wire  _T_27; 
  wire [31:0] _T_9_bits_address; 
  wire  _T_28; 
  wire  _T_29; 
  wire [31:0] _T_30; 
  wire [31:0] _T_31; 
  wire [7:0] _T_9_bits_mask; 
  wire [3:0] _T_33; 
  wire [3:0] _T_34; 
  wire  _T_37; 
  wire [9:0] _T_39; 
  wire [2:0] _T_40; 
  wire [2:0] _T_41; 
  wire  _T_42; 
  reg  _T_43; 
  reg [31:0] _RAND_1;
  wire  _T_45; 
  wire  _T_46; 
  wire  _T_47; 
  wire  _T_49; 
  wire  _T_51; 
  reg  _T_56; 
  reg [31:0] _RAND_2;
  wire  _T_57; 
  wire  _T_61; 
  wire  _T_62; 
  wire  _T_58; 
  wire  _T_60; 
  reg [31:0] _T_64_0; 
  reg [31:0] _RAND_3;
  wire [31:0] _T_65; 
  wire  _T_69; 
  dual_TLMonitor_12 dual_TLMonitor ( 
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_io_in_a_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt)
  );
  dual_Repeater_top Repeater_top ( 
    .clock(Repeater_clock),
    .reset(Repeater_reset),
    .io_repeat(Repeater_io_repeat),
    .io_enq_ready(Repeater_io_enq_ready),
    .io_enq_valid(Repeater_io_enq_valid),
    .io_enq_bits_opcode(Repeater_io_enq_bits_opcode),
    .io_enq_bits_param(Repeater_io_enq_bits_param),
    .io_enq_bits_size(Repeater_io_enq_bits_size),
    .io_enq_bits_source(Repeater_io_enq_bits_source),
    .io_enq_bits_address(Repeater_io_enq_bits_address),
    .io_enq_bits_mask(Repeater_io_enq_bits_mask),
    .io_enq_bits_data(Repeater_io_enq_bits_data),
    .io_enq_bits_corrupt(Repeater_io_enq_bits_corrupt),
    .io_deq_ready(Repeater_io_deq_ready),
    .io_deq_valid(Repeater_io_deq_valid),
    .io_deq_bits_opcode(Repeater_io_deq_bits_opcode),
    .io_deq_bits_param(Repeater_io_deq_bits_param),
    .io_deq_bits_size(Repeater_io_deq_bits_size),
    .io_deq_bits_source(Repeater_io_deq_bits_source),
    .io_deq_bits_address(Repeater_io_deq_bits_address),
    .io_deq_bits_mask(Repeater_io_deq_bits_mask),
    .io_deq_bits_data(Repeater_io_deq_bits_data),
    .io_deq_bits_corrupt(Repeater_io_deq_bits_corrupt)
  );
  assign _T_10 = Repeater_io_deq_bits_data[63:32]; 
  assign _T_11 = auto_in_a_bits_data[31:0]; 
  assign _T_12 = {_T_10,_T_11}; 
  assign _T_9_bits_opcode = Repeater_io_deq_bits_opcode; 
  assign _T_13 = _T_9_bits_opcode[2]; 
  assign _T_14 = _T_13 == 1'h0; 
  assign _T_9_bits_size = Repeater_io_deq_bits_size; 
  assign _T_16 = 10'h7 << _T_9_bits_size; 
  assign _T_17 = _T_16[2:0]; 
  assign _T_18 = ~ _T_17; 
  assign _T_19 = _T_18[2:2]; 
  assign _T_22 = _T_20 == _T_19; 
  assign _T_23 = _T_14 == 1'h0; 
  assign _T_24 = _T_22 | _T_23; 
  assign _T_9_valid = Repeater_io_deq_valid; 
  assign _T_25 = auto_out_a_ready & _T_9_valid; 
  assign _T_27 = _T_20 + 1'h1; 
  assign _T_9_bits_address = Repeater_io_deq_bits_address; 
  assign _T_28 = _T_9_bits_address[2]; 
  assign _T_29 = _T_28 | _T_20; 
  assign _T_30 = _T_12[31:0]; 
  assign _T_31 = _T_12[63:32]; 
  assign _T_9_bits_mask = Repeater_io_deq_bits_mask; 
  assign _T_33 = _T_9_bits_mask[3:0]; 
  assign _T_34 = _T_9_bits_mask[7:4]; 
  assign _T_37 = auto_out_d_bits_opcode[0]; 
  assign _T_39 = 10'h7 << auto_out_d_bits_size; 
  assign _T_40 = _T_39[2:0]; 
  assign _T_41 = ~ _T_40; 
  assign _T_42 = _T_41[2:2]; 
  assign _T_45 = _T_43 == _T_42; 
  assign _T_46 = _T_37 == 1'h0; 
  assign _T_47 = _T_45 | _T_46; 
  assign _T_49 = _T_43 & _T_42; 
  assign _T_51 = _T_49 == 1'h0; 
  assign _T_57 = auto_out_d_bits_corrupt | _T_56; 
  assign _T_61 = _T_47 == 1'h0; 
  assign _T_62 = auto_in_d_ready | _T_61; 
  assign _T_58 = _T_62 & auto_out_d_valid; 
  assign _T_60 = _T_43 + 1'h1; 
  assign _T_65 = _T_51 ? auto_out_d_bits_data : _T_64_0; 
  assign _T_69 = _T_58 & _T_61; 
  assign auto_in_a_ready = Repeater_io_enq_ready; 
  assign auto_in_d_valid = auto_out_d_valid & _T_47; 
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; 
  assign auto_in_d_bits_size = auto_out_d_bits_size; 
  assign auto_in_d_bits_source = auto_out_d_bits_source; 
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; 
  assign auto_in_d_bits_data = {auto_out_d_bits_data,_T_65}; 
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt | _T_56; 
  assign auto_out_a_valid = Repeater_io_deq_valid; 
  assign auto_out_a_bits_opcode = Repeater_io_deq_bits_opcode; 
  assign auto_out_a_bits_param = Repeater_io_deq_bits_param; 
  assign auto_out_a_bits_size = Repeater_io_deq_bits_size; 
  assign auto_out_a_bits_source = Repeater_io_deq_bits_source; 
  assign auto_out_a_bits_address = Repeater_io_deq_bits_address; 
  assign auto_out_a_bits_mask = _T_29 ? _T_34 : _T_33; 
  assign auto_out_a_bits_data = _T_29 ? _T_31 : _T_30; 
  assign auto_out_a_bits_corrupt = Repeater_io_deq_bits_corrupt; 
  assign auto_out_d_ready = auto_in_d_ready | _T_61; 
  assign TLMonitor_clock = clock; 
  assign TLMonitor_reset = reset; 
  assign TLMonitor_io_in_a_ready = Repeater_io_enq_ready; 
  assign TLMonitor_io_in_a_valid = auto_in_a_valid; 
  assign TLMonitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; 
  assign TLMonitor_io_in_a_bits_param = auto_in_a_bits_param; 
  assign TLMonitor_io_in_a_bits_size = auto_in_a_bits_size; 
  assign TLMonitor_io_in_a_bits_source = auto_in_a_bits_source; 
  assign TLMonitor_io_in_a_bits_address = auto_in_a_bits_address; 
  assign TLMonitor_io_in_a_bits_mask = auto_in_a_bits_mask; 
  assign TLMonitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; 
  assign TLMonitor_io_in_d_ready = auto_in_d_ready; 
  assign TLMonitor_io_in_d_valid = auto_out_d_valid & _T_47; 
  assign TLMonitor_io_in_d_bits_opcode = auto_out_d_bits_opcode; 
  assign TLMonitor_io_in_d_bits_param = auto_out_d_bits_param; 
  assign TLMonitor_io_in_d_bits_size = auto_out_d_bits_size; 
  assign TLMonitor_io_in_d_bits_source = auto_out_d_bits_source; 
  assign TLMonitor_io_in_d_bits_sink = auto_out_d_bits_sink; 
  assign TLMonitor_io_in_d_bits_denied = auto_out_d_bits_denied; 
  assign TLMonitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt | _T_56; 
  assign Repeater_clock = clock; 
  assign Repeater_reset = reset; 
  assign Repeater_io_repeat = _T_24 == 1'h0; 
  assign Repeater_io_enq_valid = auto_in_a_valid; 
  assign Repeater_io_enq_bits_opcode = auto_in_a_bits_opcode; 
  assign Repeater_io_enq_bits_param = auto_in_a_bits_param; 
  assign Repeater_io_enq_bits_size = auto_in_a_bits_size; 
  assign Repeater_io_enq_bits_source = auto_in_a_bits_source; 
  assign Repeater_io_enq_bits_address = auto_in_a_bits_address; 
  assign Repeater_io_enq_bits_mask = auto_in_a_bits_mask; 
  assign Repeater_io_enq_bits_data = auto_in_a_bits_data; 
  assign Repeater_io_enq_bits_corrupt = auto_in_a_bits_corrupt; 
  assign Repeater_io_deq_ready = auto_out_a_ready; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_20 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_43 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_56 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_64_0 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_20 <= 1'h0;
    end else begin
      if (_T_25) begin
        if (_T_24) begin
          _T_20 <= 1'h0;
        end else begin
          _T_20 <= _T_27;
        end
      end
    end
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      if (_T_58) begin
        if (_T_47) begin
          _T_43 <= 1'h0;
        end else begin
          _T_43 <= _T_60;
        end
      end
    end
    if (reset) begin
      _T_56 <= 1'h0;
    end else begin
      if (_T_58) begin
        if (_T_47) begin
          _T_56 <= 1'h0;
        end else begin
          _T_56 <= _T_57;
        end
      end
    end
    if (_T_69) begin
      if (_T_51) begin
        _T_64_0 <= auto_out_d_bits_data;
      end
    end
  end
endmodule
module dual_TLXbar_1( 
  input         clock, 
  input         reset, 
  output        auto_in_a_ready, 
  input         auto_in_a_valid, 
  input  [2:0]  auto_in_a_bits_opcode, 
  input  [2:0]  auto_in_a_bits_param, 
  input  [2:0]  auto_in_a_bits_size, 
  input  [2:0]  auto_in_a_bits_source, 
  input  [31:0] auto_in_a_bits_address, 
  input  [3:0]  auto_in_a_bits_mask, 
  input  [31:0] auto_in_a_bits_data, 
  input         auto_in_a_bits_corrupt, 
  input         auto_in_d_ready, 
  output        auto_in_d_valid, 
  output [2:0]  auto_in_d_bits_opcode, 
  output [1:0]  auto_in_d_bits_param, 
  output [2:0]  auto_in_d_bits_size, 
  output [2:0]  auto_in_d_bits_source, 
  output [5:0]  auto_in_d_bits_sink, 
  output        auto_in_d_bits_denied, 
  output [31:0] auto_in_d_bits_data, 
  output        auto_in_d_bits_corrupt, 
  input         auto_out_1_a_ready, 
  output        auto_out_1_a_valid, 
  output [2:0]  auto_out_1_a_bits_opcode, 
  output [2:0]  auto_out_1_a_bits_param, 
  output [2:0]  auto_out_1_a_bits_size, 
  output [2:0]  auto_out_1_a_bits_source, 
  output [28:0] auto_out_1_a_bits_address, 
  output [3:0]  auto_out_1_a_bits_mask, 
  output        auto_out_1_a_bits_corrupt, 
  output        auto_out_1_d_ready, 
  input         auto_out_1_d_valid, 
  input  [2:0]  auto_out_1_d_bits_opcode, 
  input  [1:0]  auto_out_1_d_bits_param, 
  input  [2:0]  auto_out_1_d_bits_size, 
  input  [2:0]  auto_out_1_d_bits_source, 
  input         auto_out_1_d_bits_sink, 
  input         auto_out_1_d_bits_denied, 
  input  [31:0] auto_out_1_d_bits_data, 
  input         auto_out_1_d_bits_corrupt, 
  input         auto_out_0_a_ready, 
  output        auto_out_0_a_valid, 
  output [2:0]  auto_out_0_a_bits_opcode, 
  output [2:0]  auto_out_0_a_bits_param, 
  output [2:0]  auto_out_0_a_bits_size, 
  output [2:0]  auto_out_0_a_bits_source, 
  output [31:0] auto_out_0_a_bits_address, 
  output [3:0]  auto_out_0_a_bits_mask, 
  output [31:0] auto_out_0_a_bits_data, 
  output        auto_out_0_a_bits_corrupt, 
  output        auto_out_0_d_ready, 
  input         auto_out_0_d_valid, 
  input  [2:0]  auto_out_0_d_bits_opcode, 
  input  [1:0]  auto_out_0_d_bits_param, 
  input  [2:0]  auto_out_0_d_bits_size, 
  input  [2:0]  auto_out_0_d_bits_source, 
  input  [4:0]  auto_out_0_d_bits_sink, 
  input         auto_out_0_d_bits_denied, 
  input  [31:0] auto_out_0_d_bits_data, 
  input         auto_out_0_d_bits_corrupt 
);
  wire  TLMonitor_clock; 
  wire  TLMonitor_reset; 
  wire  TLMonitor_io_in_a_ready; 
  wire  TLMonitor_io_in_a_valid; 
  wire [2:0] TLMonitor_io_in_a_bits_opcode; 
  wire [2:0] TLMonitor_io_in_a_bits_param; 
  wire [2:0] TLMonitor_io_in_a_bits_size; 
  wire [2:0] TLMonitor_io_in_a_bits_source; 
  wire [31:0] TLMonitor_io_in_a_bits_address; 
  wire [3:0] TLMonitor_io_in_a_bits_mask; 
  wire  TLMonitor_io_in_a_bits_corrupt; 
  wire  TLMonitor_io_in_d_ready; 
  wire  TLMonitor_io_in_d_valid; 
  wire [2:0] TLMonitor_io_in_d_bits_opcode; 
  wire [1:0] TLMonitor_io_in_d_bits_param; 
  wire [2:0] TLMonitor_io_in_d_bits_size; 
  wire [2:0] TLMonitor_io_in_d_bits_source; 
  wire [5:0] TLMonitor_io_in_d_bits_sink; 
  wire  TLMonitor_io_in_d_bits_denied; 
  wire  TLMonitor_io_in_d_bits_corrupt; 
  wire [31:0] _T_22; 
  wire [32:0] _T_23; 
  wire [32:0] _T_24; 
  wire [32:0] _T_25; 
  wire  _T_26; 
  wire [31:0] _T_27; 
  wire [32:0] _T_28; 
  wire [32:0] _T_29; 
  wire [32:0] _T_30; 
  wire  _T_31; 
  wire  requestAIO_0_0; 
  wire  _T_127; 
  wire [32:0] _T_34; 
  wire [32:0] _T_35; 
  wire [32:0] _T_36; 
  wire  requestAIO_0_1; 
  wire  _T_128; 
  reg [3:0] _T_161; 
  reg [31:0] _RAND_0;
  wire  _T_162; 
  wire  _T_231; 
  reg  _T_226_0; 
  reg [31:0] _RAND_1;
  wire  _T_232; 
  reg  _T_226_1; 
  reg [31:0] _RAND_2;
  wire  _T_233; 
  wire  _T_234; 
  wire  in_0_d_valid; 
  wire  _T_12; 
  wire [1:0] _T_164; 
  reg [1:0] _T_171; 
  reg [31:0] _RAND_3;
  wire [1:0] _T_172; 
  wire [1:0] _T_173; 
  wire [3:0] _T_174; 
  wire [2:0] _T_175; 
  wire [3:0] _GEN_5; 
  wire [3:0] _T_176; 
  wire [2:0] _T_178; 
  wire [3:0] _T_179; 
  wire [3:0] _GEN_6; 
  wire [3:0] _T_180; 
  wire [1:0] _T_181; 
  wire [1:0] _T_182; 
  wire [1:0] _T_183; 
  wire [1:0] _T_184; 
  wire  _T_193; 
  wire  _T_196; 
  wire  _T_227_0; 
  wire [5:0] out_0_d_bits_sink; 
  wire [50:0] _T_243; 
  wire [50:0] _T_244; 
  wire  _T_194; 
  wire  _T_197; 
  wire  _T_227_1; 
  wire [5:0] _GEN_7; 
  wire [5:0] out_1_d_bits_sink; 
  wire [50:0] _T_251; 
  wire [50:0] _T_252; 
  wire [50:0] _T_253; 
  wire [12:0] _T_111; 
  wire [5:0] _T_112; 
  wire [5:0] _T_113; 
  wire [3:0] _T_114; 
  wire  _T_115; 
  wire [3:0] beatsDO_0; 
  wire [12:0] _T_117; 
  wire [5:0] _T_118; 
  wire [5:0] _T_119; 
  wire [3:0] _T_120; 
  wire  _T_121; 
  wire [3:0] beatsDO_1; 
  wire  _T_163; 
  wire  _T_166; 
  wire  _T_168; 
  wire  _T_169; 
  wire  _T_185; 
  wire  _T_186; 
  wire [1:0] _T_187; 
  wire [2:0] _T_188; 
  wire [1:0] _T_189; 
  wire [1:0] _T_190; 
  wire  _T_200; 
  wire  _T_202; 
  wire  _T_205; 
  wire  _T_206; 
  wire  _T_209; 
  wire  _T_210; 
  wire  _T_212; 
  wire  _T_214; 
  wire  _T_216; 
  wire  _T_217; 
  wire [3:0] _T_218; 
  wire [3:0] _T_219; 
  wire [3:0] _T_220; 
  wire [3:0] _GEN_8; 
  wire [3:0] _T_223; 
  wire  _T_228_0; 
  wire  _T_228_1; 
  dual_TLMonitor_1 dual_TLMonitor ( 
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_io_in_a_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt)
  );
  assign _T_22 = auto_in_a_bits_address ^ 32'h40000000; 
  assign _T_23 = {1'b0,$signed(_T_22)}; 
  assign _T_24 = $signed(_T_23) & $signed(33'shc0000000); 
  assign _T_25 = $signed(_T_24); 
  assign _T_26 = $signed(_T_25) == $signed(33'sh0); 
  assign _T_27 = auto_in_a_bits_address ^ 32'h80000000; 
  assign _T_28 = {1'b0,$signed(_T_27)}; 
  assign _T_29 = $signed(_T_28) & $signed(33'sh80000000); 
  assign _T_30 = $signed(_T_29); 
  assign _T_31 = $signed(_T_30) == $signed(33'sh0); 
  assign requestAIO_0_0 = _T_26 | _T_31; 
  assign _T_127 = requestAIO_0_0 ? auto_out_0_a_ready : 1'h0; 
  assign _T_34 = {1'b0,$signed(auto_in_a_bits_address)}; 
  assign _T_35 = $signed(_T_34) & $signed(33'shc0000000); 
  assign _T_36 = $signed(_T_35); 
  assign requestAIO_0_1 = $signed(_T_36) == $signed(33'sh0); 
  assign _T_128 = requestAIO_0_1 ? auto_out_1_a_ready : 1'h0; 
  assign _T_162 = _T_161 == 4'h0; 
  assign _T_231 = auto_out_0_d_valid | auto_out_1_d_valid; 
  assign _T_232 = _T_226_0 ? auto_out_0_d_valid : 1'h0; 
  assign _T_233 = _T_226_1 ? auto_out_1_d_valid : 1'h0; 
  assign _T_234 = _T_232 | _T_233; 
  assign in_0_d_valid = _T_162 ? _T_231 : _T_234; 
  assign _T_12 = auto_in_d_ready & in_0_d_valid; 
  assign _T_164 = {auto_out_1_d_valid,auto_out_0_d_valid}; 
  assign _T_172 = ~ _T_171; 
  assign _T_173 = _T_164 & _T_172; 
  assign _T_174 = {_T_173,auto_out_1_d_valid,auto_out_0_d_valid}; 
  assign _T_175 = _T_174[3:1]; 
  assign _GEN_5 = {{1'd0}, _T_175}; 
  assign _T_176 = _T_174 | _GEN_5; 
  assign _T_178 = _T_176[3:1]; 
  assign _T_179 = {_T_171, 2'h0}; 
  assign _GEN_6 = {{1'd0}, _T_178}; 
  assign _T_180 = _GEN_6 | _T_179; 
  assign _T_181 = _T_180[3:2]; 
  assign _T_182 = _T_180[1:0]; 
  assign _T_183 = _T_181 & _T_182; 
  assign _T_184 = ~ _T_183; 
  assign _T_193 = _T_184[0]; 
  assign _T_196 = _T_193 & auto_out_0_d_valid; 
  assign _T_227_0 = _T_162 ? _T_196 : _T_226_0; 
  assign out_0_d_bits_sink = {{1'd0}, auto_out_0_d_bits_sink}; 
  assign _T_243 = {auto_out_0_d_bits_opcode,auto_out_0_d_bits_param,auto_out_0_d_bits_size,auto_out_0_d_bits_source,out_0_d_bits_sink,auto_out_0_d_bits_denied,auto_out_0_d_bits_data,auto_out_0_d_bits_corrupt}; 
  assign _T_244 = _T_227_0 ? _T_243 : 51'h0; 
  assign _T_194 = _T_184[1]; 
  assign _T_197 = _T_194 & auto_out_1_d_valid; 
  assign _T_227_1 = _T_162 ? _T_197 : _T_226_1; 
  assign _GEN_7 = {{5'd0}, auto_out_1_d_bits_sink}; 
  assign out_1_d_bits_sink = _GEN_7 | 6'h20; 
  assign _T_251 = {auto_out_1_d_bits_opcode,auto_out_1_d_bits_param,auto_out_1_d_bits_size,auto_out_1_d_bits_source,out_1_d_bits_sink,auto_out_1_d_bits_denied,auto_out_1_d_bits_data,auto_out_1_d_bits_corrupt}; 
  assign _T_252 = _T_227_1 ? _T_251 : 51'h0; 
  assign _T_253 = _T_244 | _T_252; 
  assign _T_111 = 13'h3f << auto_out_0_d_bits_size; 
  assign _T_112 = _T_111[5:0]; 
  assign _T_113 = ~ _T_112; 
  assign _T_114 = _T_113[5:2]; 
  assign _T_115 = auto_out_0_d_bits_opcode[0]; 
  assign beatsDO_0 = _T_115 ? _T_114 : 4'h0; 
  assign _T_117 = 13'h3f << auto_out_1_d_bits_size; 
  assign _T_118 = _T_117[5:0]; 
  assign _T_119 = ~ _T_118; 
  assign _T_120 = _T_119[5:2]; 
  assign _T_121 = auto_out_1_d_bits_opcode[0]; 
  assign beatsDO_1 = _T_121 ? _T_120 : 4'h0; 
  assign _T_163 = _T_162 & auto_in_d_ready; 
  assign _T_166 = _T_164 == _T_164; 
  assign _T_168 = _T_166 | reset; 
  assign _T_169 = _T_168 == 1'h0; 
  assign _T_185 = _T_164 != 2'h0; 
  assign _T_186 = _T_163 & _T_185; 
  assign _T_187 = _T_184 & _T_164; 
  assign _T_188 = {_T_187, 1'h0}; 
  assign _T_189 = _T_188[1:0]; 
  assign _T_190 = _T_187 | _T_189; 
  assign _T_200 = _T_196 | _T_197; 
  assign _T_202 = _T_196 == 1'h0; 
  assign _T_205 = _T_197 == 1'h0; 
  assign _T_206 = _T_202 | _T_205; 
  assign _T_209 = _T_206 | reset; 
  assign _T_210 = _T_209 == 1'h0; 
  assign _T_212 = _T_231 == 1'h0; 
  assign _T_214 = _T_212 | _T_200; 
  assign _T_216 = _T_214 | reset; 
  assign _T_217 = _T_216 == 1'h0; 
  assign _T_218 = _T_196 ? beatsDO_0 : 4'h0; 
  assign _T_219 = _T_197 ? beatsDO_1 : 4'h0; 
  assign _T_220 = _T_218 | _T_219; 
  assign _GEN_8 = {{3'd0}, _T_12}; 
  assign _T_223 = _T_161 - _GEN_8; 
  assign _T_228_0 = _T_162 ? _T_193 : _T_226_0; 
  assign _T_228_1 = _T_162 ? _T_194 : _T_226_1; 
  assign auto_in_a_ready = _T_127 | _T_128; 
  assign auto_in_d_valid = _T_162 ? _T_231 : _T_234; 
  assign auto_in_d_bits_opcode = _T_253[50:48]; 
  assign auto_in_d_bits_param = _T_253[47:46]; 
  assign auto_in_d_bits_size = _T_253[45:43]; 
  assign auto_in_d_bits_source = _T_253[42:40]; 
  assign auto_in_d_bits_sink = _T_253[39:34]; 
  assign auto_in_d_bits_denied = _T_253[33]; 
  assign auto_in_d_bits_data = _T_253[32:1]; 
  assign auto_in_d_bits_corrupt = _T_253[0]; 
  assign auto_out_1_a_valid = auto_in_a_valid & requestAIO_0_1; 
  assign auto_out_1_a_bits_opcode = auto_in_a_bits_opcode; 
  assign auto_out_1_a_bits_param = auto_in_a_bits_param; 
  assign auto_out_1_a_bits_size = auto_in_a_bits_size; 
  assign auto_out_1_a_bits_source = auto_in_a_bits_source; 
  assign auto_out_1_a_bits_address = auto_in_a_bits_address[28:0]; 
  assign auto_out_1_a_bits_mask = auto_in_a_bits_mask; 
  assign auto_out_1_a_bits_corrupt = auto_in_a_bits_corrupt; 
  assign auto_out_1_d_ready = auto_in_d_ready & _T_228_1; 
  assign auto_out_0_a_valid = auto_in_a_valid & requestAIO_0_0; 
  assign auto_out_0_a_bits_opcode = auto_in_a_bits_opcode; 
  assign auto_out_0_a_bits_param = auto_in_a_bits_param; 
  assign auto_out_0_a_bits_size = auto_in_a_bits_size; 
  assign auto_out_0_a_bits_source = auto_in_a_bits_source; 
  assign auto_out_0_a_bits_address = auto_in_a_bits_address; 
  assign auto_out_0_a_bits_mask = auto_in_a_bits_mask; 
  assign auto_out_0_a_bits_data = auto_in_a_bits_data; 
  assign auto_out_0_a_bits_corrupt = auto_in_a_bits_corrupt; 
  assign auto_out_0_d_ready = auto_in_d_ready & _T_228_0; 
  assign TLMonitor_clock = clock; 
  assign TLMonitor_reset = reset; 
  assign TLMonitor_io_in_a_ready = _T_127 | _T_128; 
  assign TLMonitor_io_in_a_valid = auto_in_a_valid; 
  assign TLMonitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; 
  assign TLMonitor_io_in_a_bits_param = auto_in_a_bits_param; 
  assign TLMonitor_io_in_a_bits_size = auto_in_a_bits_size; 
  assign TLMonitor_io_in_a_bits_source = auto_in_a_bits_source; 
  assign TLMonitor_io_in_a_bits_address = auto_in_a_bits_address; 
  assign TLMonitor_io_in_a_bits_mask = auto_in_a_bits_mask; 
  assign TLMonitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; 
  assign TLMonitor_io_in_d_ready = auto_in_d_ready; 
  assign TLMonitor_io_in_d_valid = _T_162 ? _T_231 : _T_234; 
  assign TLMonitor_io_in_d_bits_opcode = _T_253[50:48]; 
  assign TLMonitor_io_in_d_bits_param = _T_253[47:46]; 
  assign TLMonitor_io_in_d_bits_size = _T_253[45:43]; 
  assign TLMonitor_io_in_d_bits_source = _T_253[42:40]; 
  assign TLMonitor_io_in_d_bits_sink = _T_253[39:34]; 
  assign TLMonitor_io_in_d_bits_denied = _T_253[33]; 
  assign TLMonitor_io_in_d_bits_corrupt = _T_253[0]; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_161 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_226_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_226_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_171 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_161 <= 4'h0;
    end else begin
      if (_T_163) begin
        _T_161 <= _T_220;
      end else begin
        _T_161 <= _T_223;
      end
    end
    if (reset) begin
      _T_226_0 <= 1'h0;
    end else begin
      if (_T_162) begin
        _T_226_0 <= _T_196;
      end
    end
    if (reset) begin
      _T_226_1 <= 1'h0;
    end else begin
      if (_T_162) begin
        _T_226_1 <= _T_197;
      end
    end
    if (reset) begin
      _T_171 <= 2'h3;
    end else begin
      if (_T_186) begin
        _T_171 <= _T_190;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_169) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_169) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_210) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_210) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_217) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:70 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_217) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TLXbar( 
  input         clock, 
  input         reset, 
  output        auto_in_a_ready, 
  input         auto_in_a_valid, 
  input  [2:0]  auto_in_a_bits_opcode, 
  input  [2:0]  auto_in_a_bits_param, 
  input  [3:0]  auto_in_a_bits_size, 
  input  [6:0]  auto_in_a_bits_source, 
  input  [31:0] auto_in_a_bits_address, 
  input  [7:0]  auto_in_a_bits_mask, 
  input  [63:0] auto_in_a_bits_data, 
  input         auto_in_a_bits_corrupt, 
  output        auto_in_c_ready, 
  input         auto_in_c_valid, 
  input  [2:0]  auto_in_c_bits_opcode, 
  input  [2:0]  auto_in_c_bits_param, 
  input  [3:0]  auto_in_c_bits_size, 
  input  [6:0]  auto_in_c_bits_source, 
  input  [31:0] auto_in_c_bits_address, 
  input         auto_in_c_bits_corrupt, 
  input         auto_in_d_ready, 
  output        auto_in_d_valid, 
  output [2:0]  auto_in_d_bits_opcode, 
  output [1:0]  auto_in_d_bits_param, 
  output [3:0]  auto_in_d_bits_size, 
  output [6:0]  auto_in_d_bits_source, 
  output        auto_in_d_bits_sink, 
  output        auto_in_d_bits_denied, 
  output [63:0] auto_in_d_bits_data, 
  output        auto_in_d_bits_corrupt, 
  output        auto_in_e_ready, 
  input         auto_in_e_valid, 
  input         auto_in_e_bits_sink, 
  input         auto_out_2_a_ready, 
  output        auto_out_2_a_valid, 
  output [2:0]  auto_out_2_a_bits_opcode, 
  output [2:0]  auto_out_2_a_bits_param, 
  output [2:0]  auto_out_2_a_bits_size, 
  output [6:0]  auto_out_2_a_bits_source, 
  output [28:0] auto_out_2_a_bits_address, 
  output [7:0]  auto_out_2_a_bits_mask, 
  output        auto_out_2_a_bits_corrupt, 
  input         auto_out_2_c_ready, 
  output        auto_out_2_c_valid, 
  output [2:0]  auto_out_2_c_bits_opcode, 
  output [2:0]  auto_out_2_c_bits_param, 
  output [2:0]  auto_out_2_c_bits_size, 
  output [6:0]  auto_out_2_c_bits_source, 
  output [28:0] auto_out_2_c_bits_address, 
  output        auto_out_2_c_bits_corrupt, 
  output        auto_out_2_d_ready, 
  input         auto_out_2_d_valid, 
  input  [2:0]  auto_out_2_d_bits_opcode, 
  input  [1:0]  auto_out_2_d_bits_param, 
  input  [2:0]  auto_out_2_d_bits_size, 
  input  [6:0]  auto_out_2_d_bits_source, 
  input         auto_out_2_d_bits_sink, 
  input         auto_out_2_d_bits_denied, 
  input  [63:0] auto_out_2_d_bits_data, 
  input         auto_out_2_d_bits_corrupt, 
  output        auto_out_2_e_valid, 
  input         auto_out_1_a_ready, 
  output        auto_out_1_a_valid, 
  output [2:0]  auto_out_1_a_bits_opcode, 
  output [2:0]  auto_out_1_a_bits_param, 
  output [3:0]  auto_out_1_a_bits_size, 
  output [6:0]  auto_out_1_a_bits_source, 
  output [30:0] auto_out_1_a_bits_address, 
  output [7:0]  auto_out_1_a_bits_mask, 
  output [63:0] auto_out_1_a_bits_data, 
  output        auto_out_1_a_bits_corrupt, 
  output        auto_out_1_d_ready, 
  input         auto_out_1_d_valid, 
  input  [2:0]  auto_out_1_d_bits_opcode, 
  input  [3:0]  auto_out_1_d_bits_size, 
  input  [6:0]  auto_out_1_d_bits_source, 
  input         auto_out_1_d_bits_denied, 
  input  [63:0] auto_out_1_d_bits_data, 
  input         auto_out_1_d_bits_corrupt, 
  input         auto_out_0_a_ready, 
  output        auto_out_0_a_valid, 
  output [2:0]  auto_out_0_a_bits_opcode, 
  output [2:0]  auto_out_0_a_bits_param, 
  output [2:0]  auto_out_0_a_bits_size, 
  output [6:0]  auto_out_0_a_bits_source, 
  output [31:0] auto_out_0_a_bits_address, 
  output [7:0]  auto_out_0_a_bits_mask, 
  output [63:0] auto_out_0_a_bits_data, 
  output        auto_out_0_a_bits_corrupt, 
  output        auto_out_0_d_ready, 
  input         auto_out_0_d_valid, 
  input  [2:0]  auto_out_0_d_bits_opcode, 
  input  [2:0]  auto_out_0_d_bits_size, 
  input  [6:0]  auto_out_0_d_bits_source, 
  input         auto_out_0_d_bits_denied, 
  input  [63:0] auto_out_0_d_bits_data, 
  input         auto_out_0_d_bits_corrupt 
);
  wire  TLMonitor_clock; 
  wire  TLMonitor_reset; 
  wire  TLMonitor_io_in_a_ready; 
  wire  TLMonitor_io_in_a_valid; 
  wire [2:0] TLMonitor_io_in_a_bits_opcode; 
  wire [2:0] TLMonitor_io_in_a_bits_param; 
  wire [3:0] TLMonitor_io_in_a_bits_size; 
  wire [6:0] TLMonitor_io_in_a_bits_source; 
  wire [31:0] TLMonitor_io_in_a_bits_address; 
  wire [7:0] TLMonitor_io_in_a_bits_mask; 
  wire  TLMonitor_io_in_a_bits_corrupt; 
  wire  TLMonitor_io_in_c_ready; 
  wire  TLMonitor_io_in_c_valid; 
  wire [2:0] TLMonitor_io_in_c_bits_opcode; 
  wire [2:0] TLMonitor_io_in_c_bits_param; 
  wire [3:0] TLMonitor_io_in_c_bits_size; 
  wire [6:0] TLMonitor_io_in_c_bits_source; 
  wire [31:0] TLMonitor_io_in_c_bits_address; 
  wire  TLMonitor_io_in_c_bits_corrupt; 
  wire  TLMonitor_io_in_d_ready; 
  wire  TLMonitor_io_in_d_valid; 
  wire [2:0] TLMonitor_io_in_d_bits_opcode; 
  wire [1:0] TLMonitor_io_in_d_bits_param; 
  wire [3:0] TLMonitor_io_in_d_bits_size; 
  wire [6:0] TLMonitor_io_in_d_bits_source; 
  wire  TLMonitor_io_in_d_bits_sink; 
  wire  TLMonitor_io_in_d_bits_denied; 
  wire  TLMonitor_io_in_d_bits_corrupt; 
  wire  TLMonitor_io_in_e_ready; 
  wire  TLMonitor_io_in_e_valid; 
  wire  TLMonitor_io_in_e_bits_sink; 
  wire [31:0] _T_25; 
  wire [32:0] _T_26; 
  wire [32:0] _T_27; 
  wire [32:0] _T_28; 
  wire  requestAIO_0_0; 
  wire  _T_156; 
  wire [31:0] _T_30; 
  wire [32:0] _T_31; 
  wire [32:0] _T_32; 
  wire [32:0] _T_33; 
  wire  requestAIO_0_1; 
  wire  _T_157; 
  wire  _T_159; 
  wire [32:0] _T_36; 
  wire [32:0] _T_37; 
  wire [32:0] _T_38; 
  wire  requestAIO_0_2; 
  wire  _T_158; 
  reg [4:0] _T_206; 
  reg [31:0] _RAND_0;
  wire  _T_207; 
  wire  _T_294; 
  wire  _T_295; 
  reg  _T_288_0; 
  reg [31:0] _RAND_1;
  wire  _T_296; 
  reg  _T_288_1; 
  reg [31:0] _RAND_2;
  wire  _T_297; 
  wire  _T_299; 
  reg  _T_288_2; 
  reg [31:0] _RAND_3;
  wire  _T_298; 
  wire  _T_300; 
  wire  in_0_d_valid; 
  wire  _T_12; 
  wire [2:0] _T_210; 
  reg [2:0] _T_217; 
  reg [31:0] _RAND_4;
  wire [2:0] _T_218; 
  wire [2:0] _T_219; 
  wire [5:0] _T_220; 
  wire [4:0] _T_221; 
  wire [5:0] _GEN_5; 
  wire [5:0] _T_222; 
  wire [3:0] _T_223; 
  wire [5:0] _GEN_6; 
  wire [5:0] _T_224; 
  wire [4:0] _T_226; 
  wire [5:0] _T_227; 
  wire [5:0] _GEN_7; 
  wire [5:0] _T_228; 
  wire [2:0] _T_229; 
  wire [2:0] _T_230; 
  wire [2:0] _T_231; 
  wire [2:0] _T_232; 
  wire  _T_244; 
  wire  _T_248; 
  wire  _T_289_0; 
  wire [3:0] out_0_d_bits_size; 
  wire [82:0] _T_309; 
  wire [82:0] _T_310; 
  wire  _T_245; 
  wire  _T_249; 
  wire  _T_289_1; 
  wire [82:0] _T_317; 
  wire [82:0] _T_318; 
  wire [82:0] _T_327; 
  wire  _T_246; 
  wire  _T_250; 
  wire  _T_289_2; 
  wire [3:0] out_2_d_bits_size; 
  wire [82:0] _T_325; 
  wire [82:0] _T_326; 
  wire [82:0] _T_328; 
  wire  requestEIO_0_2; 
  wire [20:0] _T_132; 
  wire [5:0] _T_133; 
  wire [5:0] _T_134; 
  wire [2:0] _T_135; 
  wire  _T_136; 
  wire [2:0] beatsDO_0; 
  wire [22:0] _T_138; 
  wire [7:0] _T_139; 
  wire [7:0] _T_140; 
  wire [4:0] _T_141; 
  wire  _T_142; 
  wire [4:0] beatsDO_1; 
  wire [20:0] _T_144; 
  wire [5:0] _T_145; 
  wire [5:0] _T_146; 
  wire [2:0] _T_147; 
  wire  _T_148; 
  wire [2:0] beatsDO_2; 
  wire  _T_208; 
  wire  _T_212; 
  wire  _T_214; 
  wire  _T_215; 
  wire  _T_233; 
  wire  _T_234; 
  wire [2:0] _T_235; 
  wire [3:0] _T_236; 
  wire [2:0] _T_237; 
  wire [2:0] _T_238; 
  wire [4:0] _T_239; 
  wire [2:0] _T_240; 
  wire [2:0] _T_241; 
  wire  _T_253; 
  wire  _T_254; 
  wire  _T_256; 
  wire  _T_259; 
  wire  _T_260; 
  wire  _T_261; 
  wire  _T_262; 
  wire  _T_263; 
  wire  _T_265; 
  wire  _T_267; 
  wire  _T_268; 
  wire  _T_271; 
  wire  _T_274; 
  wire  _T_276; 
  wire  _T_277; 
  wire [2:0] _T_278; 
  wire [4:0] _T_279; 
  wire [2:0] _T_280; 
  wire [4:0] _GEN_8; 
  wire [4:0] _T_281; 
  wire [4:0] _GEN_9; 
  wire [4:0] _T_282; 
  wire [4:0] _GEN_10; 
  wire [4:0] _T_285; 
  wire  _T_290_0; 
  wire  _T_290_1; 
  wire  _T_290_2; 
  dual_TLMonitor TLMonitor ( 
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_io_in_a_bits_corrupt),
    .io_in_c_ready(TLMonitor_io_in_c_ready),
    .io_in_c_valid(TLMonitor_io_in_c_valid),
    .io_in_c_bits_opcode(TLMonitor_io_in_c_bits_opcode),
    .io_in_c_bits_param(TLMonitor_io_in_c_bits_param),
    .io_in_c_bits_size(TLMonitor_io_in_c_bits_size),
    .io_in_c_bits_source(TLMonitor_io_in_c_bits_source),
    .io_in_c_bits_address(TLMonitor_io_in_c_bits_address),
    .io_in_c_bits_corrupt(TLMonitor_io_in_c_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(TLMonitor_io_in_d_bits_param),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source),
    .io_in_d_bits_sink(TLMonitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(TLMonitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(TLMonitor_io_in_d_bits_corrupt),
    .io_in_e_ready(TLMonitor_io_in_e_ready),
    .io_in_e_valid(TLMonitor_io_in_e_valid),
    .io_in_e_bits_sink(TLMonitor_io_in_e_bits_sink)
  );
  assign _T_25 = auto_in_a_bits_address ^ 32'h80000000; 
  assign _T_26 = {1'b0,$signed(_T_25)}; 
  assign _T_27 = $signed(_T_26) & $signed(33'sh80000000); 
  assign _T_28 = $signed(_T_27); 
  assign requestAIO_0_0 = $signed(_T_28) == $signed(33'sh0); 
  assign _T_156 = requestAIO_0_0 ? auto_out_0_a_ready : 1'h0; 
  assign _T_30 = auto_in_a_bits_address ^ 32'h40000000; 
  assign _T_31 = {1'b0,$signed(_T_30)}; 
  assign _T_32 = $signed(_T_31) & $signed(33'shc0000000); 
  assign _T_33 = $signed(_T_32); 
  assign requestAIO_0_1 = $signed(_T_33) == $signed(33'sh0); 
  assign _T_157 = requestAIO_0_1 ? auto_out_1_a_ready : 1'h0; 
  assign _T_159 = _T_156 | _T_157; 
  assign _T_36 = {1'b0,$signed(auto_in_a_bits_address)}; 
  assign _T_37 = $signed(_T_36) & $signed(33'shc0000000); 
  assign _T_38 = $signed(_T_37); 
  assign requestAIO_0_2 = $signed(_T_38) == $signed(33'sh0); 
  assign _T_158 = requestAIO_0_2 ? auto_out_2_a_ready : 1'h0; 
  assign _T_207 = _T_206 == 5'h0; 
  assign _T_294 = auto_out_0_d_valid | auto_out_1_d_valid; 
  assign _T_295 = _T_294 | auto_out_2_d_valid; 
  assign _T_296 = _T_288_0 ? auto_out_0_d_valid : 1'h0; 
  assign _T_297 = _T_288_1 ? auto_out_1_d_valid : 1'h0; 
  assign _T_299 = _T_296 | _T_297; 
  assign _T_298 = _T_288_2 ? auto_out_2_d_valid : 1'h0; 
  assign _T_300 = _T_299 | _T_298; 
  assign in_0_d_valid = _T_207 ? _T_295 : _T_300; 
  assign _T_12 = auto_in_d_ready & in_0_d_valid; 
  assign _T_210 = {auto_out_2_d_valid,auto_out_1_d_valid,auto_out_0_d_valid}; 
  assign _T_218 = ~ _T_217; 
  assign _T_219 = _T_210 & _T_218; 
  assign _T_220 = {_T_219,auto_out_2_d_valid,auto_out_1_d_valid,auto_out_0_d_valid}; 
  assign _T_221 = _T_220[5:1]; 
  assign _GEN_5 = {{1'd0}, _T_221}; 
  assign _T_222 = _T_220 | _GEN_5; 
  assign _T_223 = _T_222[5:2]; 
  assign _GEN_6 = {{2'd0}, _T_223}; 
  assign _T_224 = _T_222 | _GEN_6; 
  assign _T_226 = _T_224[5:1]; 
  assign _T_227 = {_T_217, 3'h0}; 
  assign _GEN_7 = {{1'd0}, _T_226}; 
  assign _T_228 = _GEN_7 | _T_227; 
  assign _T_229 = _T_228[5:3]; 
  assign _T_230 = _T_228[2:0]; 
  assign _T_231 = _T_229 & _T_230; 
  assign _T_232 = ~ _T_231; 
  assign _T_244 = _T_232[0]; 
  assign _T_248 = _T_244 & auto_out_0_d_valid; 
  assign _T_289_0 = _T_207 ? _T_248 : _T_288_0; 
  assign out_0_d_bits_size = {{1'd0}, auto_out_0_d_bits_size}; 
  assign _T_309 = {auto_out_0_d_bits_opcode,2'h0,out_0_d_bits_size,auto_out_0_d_bits_source,1'h0,auto_out_0_d_bits_denied,auto_out_0_d_bits_data,auto_out_0_d_bits_corrupt}; 
  assign _T_310 = _T_289_0 ? _T_309 : 83'h0; 
  assign _T_245 = _T_232[1]; 
  assign _T_249 = _T_245 & auto_out_1_d_valid; 
  assign _T_289_1 = _T_207 ? _T_249 : _T_288_1; 
  assign _T_317 = {auto_out_1_d_bits_opcode,2'h0,auto_out_1_d_bits_size,auto_out_1_d_bits_source,1'h0,auto_out_1_d_bits_denied,auto_out_1_d_bits_data,auto_out_1_d_bits_corrupt}; 
  assign _T_318 = _T_289_1 ? _T_317 : 83'h0; 
  assign _T_327 = _T_310 | _T_318; 
  assign _T_246 = _T_232[2]; 
  assign _T_250 = _T_246 & auto_out_2_d_valid; 
  assign _T_289_2 = _T_207 ? _T_250 : _T_288_2; 
  assign out_2_d_bits_size = {{1'd0}, auto_out_2_d_bits_size}; 
  assign _T_325 = {auto_out_2_d_bits_opcode,auto_out_2_d_bits_param,out_2_d_bits_size,auto_out_2_d_bits_source,auto_out_2_d_bits_sink,auto_out_2_d_bits_denied,auto_out_2_d_bits_data,auto_out_2_d_bits_corrupt}; 
  assign _T_326 = _T_289_2 ? _T_325 : 83'h0; 
  assign _T_328 = _T_327 | _T_326; 
  assign requestEIO_0_2 = auto_in_e_bits_sink == 1'h0; 
  assign _T_132 = 21'h3f << out_0_d_bits_size; 
  assign _T_133 = _T_132[5:0]; 
  assign _T_134 = ~ _T_133; 
  assign _T_135 = _T_134[5:3]; 
  assign _T_136 = auto_out_0_d_bits_opcode[0]; 
  assign beatsDO_0 = _T_136 ? _T_135 : 3'h0; 
  assign _T_138 = 23'hff << auto_out_1_d_bits_size; 
  assign _T_139 = _T_138[7:0]; 
  assign _T_140 = ~ _T_139; 
  assign _T_141 = _T_140[7:3]; 
  assign _T_142 = auto_out_1_d_bits_opcode[0]; 
  assign beatsDO_1 = _T_142 ? _T_141 : 5'h0; 
  assign _T_144 = 21'h3f << out_2_d_bits_size; 
  assign _T_145 = _T_144[5:0]; 
  assign _T_146 = ~ _T_145; 
  assign _T_147 = _T_146[5:3]; 
  assign _T_148 = auto_out_2_d_bits_opcode[0]; 
  assign beatsDO_2 = _T_148 ? _T_147 : 3'h0; 
  assign _T_208 = _T_207 & auto_in_d_ready; 
  assign _T_212 = _T_210 == _T_210; 
  assign _T_214 = _T_212 | reset; 
  assign _T_215 = _T_214 == 1'h0; 
  assign _T_233 = _T_210 != 3'h0; 
  assign _T_234 = _T_208 & _T_233; 
  assign _T_235 = _T_232 & _T_210; 
  assign _T_236 = {_T_235, 1'h0}; 
  assign _T_237 = _T_236[2:0]; 
  assign _T_238 = _T_235 | _T_237; 
  assign _T_239 = {_T_238, 2'h0}; 
  assign _T_240 = _T_239[2:0]; 
  assign _T_241 = _T_238 | _T_240; 
  assign _T_253 = _T_248 | _T_249; 
  assign _T_254 = _T_253 | _T_250; 
  assign _T_256 = _T_248 == 1'h0; 
  assign _T_259 = _T_249 == 1'h0; 
  assign _T_260 = _T_256 | _T_259; 
  assign _T_261 = _T_253 == 1'h0; 
  assign _T_262 = _T_250 == 1'h0; 
  assign _T_263 = _T_261 | _T_262; 
  assign _T_265 = _T_260 & _T_263; 
  assign _T_267 = _T_265 | reset; 
  assign _T_268 = _T_267 == 1'h0; 
  assign _T_271 = _T_295 == 1'h0; 
  assign _T_274 = _T_271 | _T_254; 
  assign _T_276 = _T_274 | reset; 
  assign _T_277 = _T_276 == 1'h0; 
  assign _T_278 = _T_248 ? beatsDO_0 : 3'h0; 
  assign _T_279 = _T_249 ? beatsDO_1 : 5'h0; 
  assign _T_280 = _T_250 ? beatsDO_2 : 3'h0; 
  assign _GEN_8 = {{2'd0}, _T_278}; 
  assign _T_281 = _GEN_8 | _T_279; 
  assign _GEN_9 = {{2'd0}, _T_280}; 
  assign _T_282 = _T_281 | _GEN_9; 
  assign _GEN_10 = {{4'd0}, _T_12}; 
  assign _T_285 = _T_206 - _GEN_10; 
  assign _T_290_0 = _T_207 ? _T_244 : _T_288_0; 
  assign _T_290_1 = _T_207 ? _T_245 : _T_288_1; 
  assign _T_290_2 = _T_207 ? _T_246 : _T_288_2; 
  assign auto_in_a_ready = _T_159 | _T_158; 
  assign auto_in_c_ready = auto_out_2_c_ready; 
  assign auto_in_d_valid = _T_207 ? _T_295 : _T_300; 
  assign auto_in_d_bits_opcode = _T_328[82:80]; 
  assign auto_in_d_bits_param = _T_328[79:78]; 
  assign auto_in_d_bits_size = _T_328[77:74]; 
  assign auto_in_d_bits_source = _T_328[73:67]; 
  assign auto_in_d_bits_sink = _T_328[66]; 
  assign auto_in_d_bits_denied = _T_328[65]; 
  assign auto_in_d_bits_data = _T_328[64:1]; 
  assign auto_in_d_bits_corrupt = _T_328[0]; 
  assign auto_in_e_ready = auto_in_e_bits_sink == 1'h0; 
  assign auto_out_2_a_valid = auto_in_a_valid & requestAIO_0_2; 
  assign auto_out_2_a_bits_opcode = auto_in_a_bits_opcode; 
  assign auto_out_2_a_bits_param = auto_in_a_bits_param; 
  assign auto_out_2_a_bits_size = auto_in_a_bits_size[2:0]; 
  assign auto_out_2_a_bits_source = auto_in_a_bits_source; 
  assign auto_out_2_a_bits_address = auto_in_a_bits_address[28:0]; 
  assign auto_out_2_a_bits_mask = auto_in_a_bits_mask; 
  assign auto_out_2_a_bits_corrupt = auto_in_a_bits_corrupt; 
  assign auto_out_2_c_valid = auto_in_c_valid; 
  assign auto_out_2_c_bits_opcode = auto_in_c_bits_opcode; 
  assign auto_out_2_c_bits_param = auto_in_c_bits_param; 
  assign auto_out_2_c_bits_size = auto_in_c_bits_size[2:0]; 
  assign auto_out_2_c_bits_source = auto_in_c_bits_source; 
  assign auto_out_2_c_bits_address = auto_in_c_bits_address[28:0]; 
  assign auto_out_2_c_bits_corrupt = auto_in_c_bits_corrupt; 
  assign auto_out_2_d_ready = auto_in_d_ready & _T_290_2; 
  assign auto_out_2_e_valid = auto_in_e_valid & requestEIO_0_2; 
  assign auto_out_1_a_valid = auto_in_a_valid & requestAIO_0_1; 
  assign auto_out_1_a_bits_opcode = auto_in_a_bits_opcode; 
  assign auto_out_1_a_bits_param = auto_in_a_bits_param; 
  assign auto_out_1_a_bits_size = auto_in_a_bits_size; 
  assign auto_out_1_a_bits_source = auto_in_a_bits_source; 
  assign auto_out_1_a_bits_address = auto_in_a_bits_address[30:0]; 
  assign auto_out_1_a_bits_mask = auto_in_a_bits_mask; 
  assign auto_out_1_a_bits_data = auto_in_a_bits_data; 
  assign auto_out_1_a_bits_corrupt = auto_in_a_bits_corrupt; 
  assign auto_out_1_d_ready = auto_in_d_ready & _T_290_1; 
  assign auto_out_0_a_valid = auto_in_a_valid & requestAIO_0_0; 
  assign auto_out_0_a_bits_opcode = auto_in_a_bits_opcode; 
  assign auto_out_0_a_bits_param = auto_in_a_bits_param; 
  assign auto_out_0_a_bits_size = auto_in_a_bits_size[2:0]; 
  assign auto_out_0_a_bits_source = auto_in_a_bits_source; 
  assign auto_out_0_a_bits_address = auto_in_a_bits_address; 
  assign auto_out_0_a_bits_mask = auto_in_a_bits_mask; 
  assign auto_out_0_a_bits_data = auto_in_a_bits_data; 
  assign auto_out_0_a_bits_corrupt = auto_in_a_bits_corrupt; 
  assign auto_out_0_d_ready = auto_in_d_ready & _T_290_0; 
  assign TLMonitor_clock = clock; 
  assign TLMonitor_reset = reset; 
  assign TLMonitor_io_in_a_ready = _T_159 | _T_158; 
  assign TLMonitor_io_in_a_valid = auto_in_a_valid; 
  assign TLMonitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; 
  assign TLMonitor_io_in_a_bits_param = auto_in_a_bits_param; 
  assign TLMonitor_io_in_a_bits_size = auto_in_a_bits_size; 
  assign TLMonitor_io_in_a_bits_source = auto_in_a_bits_source; 
  assign TLMonitor_io_in_a_bits_address = auto_in_a_bits_address; 
  assign TLMonitor_io_in_a_bits_mask = auto_in_a_bits_mask; 
  assign TLMonitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; 
  assign TLMonitor_io_in_c_ready = auto_out_2_c_ready; 
  assign TLMonitor_io_in_c_valid = auto_in_c_valid; 
  assign TLMonitor_io_in_c_bits_opcode = auto_in_c_bits_opcode; 
  assign TLMonitor_io_in_c_bits_param = auto_in_c_bits_param; 
  assign TLMonitor_io_in_c_bits_size = auto_in_c_bits_size; 
  assign TLMonitor_io_in_c_bits_source = auto_in_c_bits_source; 
  assign TLMonitor_io_in_c_bits_address = auto_in_c_bits_address; 
  assign TLMonitor_io_in_c_bits_corrupt = auto_in_c_bits_corrupt; 
  assign TLMonitor_io_in_d_ready = auto_in_d_ready; 
  assign TLMonitor_io_in_d_valid = _T_207 ? _T_295 : _T_300; 
  assign TLMonitor_io_in_d_bits_opcode = _T_328[82:80]; 
  assign TLMonitor_io_in_d_bits_param = _T_328[79:78]; 
  assign TLMonitor_io_in_d_bits_size = _T_328[77:74]; 
  assign TLMonitor_io_in_d_bits_source = _T_328[73:67]; 
  assign TLMonitor_io_in_d_bits_sink = _T_328[66]; 
  assign TLMonitor_io_in_d_bits_denied = _T_328[65]; 
  assign TLMonitor_io_in_d_bits_corrupt = _T_328[0]; 
  assign TLMonitor_io_in_e_ready = auto_in_e_bits_sink == 1'h0; 
  assign TLMonitor_io_in_e_valid = auto_in_e_valid; 
  assign TLMonitor_io_in_e_bits_sink = auto_in_e_bits_sink; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_206 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_288_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_288_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_288_2 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_217 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_206 <= 5'h0;
    end else begin
      if (_T_208) begin
        _T_206 <= _T_282;
      end else begin
        _T_206 <= _T_285;
      end
    end
    if (reset) begin
      _T_288_0 <= 1'h0;
    end else begin
      if (_T_207) begin
        _T_288_0 <= _T_248;
      end
    end
    if (reset) begin
      _T_288_1 <= 1'h0;
    end else begin
      if (_T_207) begin
        _T_288_1 <= _T_249;
      end
    end
    if (reset) begin
      _T_288_2 <= 1'h0;
    end else begin
      if (_T_207) begin
        _T_288_2 <= _T_250;
      end
    end
    if (reset) begin
      _T_217 <= 3'h7;
    end else begin
      if (_T_234) begin
        _T_217 <= _T_241;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_215) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_215) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_268) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_268) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_277) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:70 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_277) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module dual_TX( 
  input         clock, 
  input         reset, 
  output        io_c2b_clk, 
  output        io_c2b_rst, 
  output        io_c2b_send, 
  output [31:0] io_c2b_data, 
  output        io_sa_ready, 
  input         io_sa_valid, 
  input  [31:0] io_sa_bits_data, 
  input         io_sa_bits_last, 
  input  [12:0] io_sa_bits_beats, 
  output        io_sb_ready, 
  input  [31:0] io_sb_bits_data, 
  input         io_sb_bits_last, 
  output        io_sc_ready, 
  input  [31:0] io_sc_bits_data, 
  input         io_sc_bits_last, 
  output        io_sd_ready, 
  input         io_sd_valid, 
  input  [31:0] io_sd_bits_data, 
  input         io_sd_bits_last, 
  input  [12:0] io_sd_bits_beats, 
  input  [31:0] io_se_bits_data, 
  input  [19:0] io_rxc_mem_0_a, 
  input  [19:0] io_rxc_mem_0_b, 
  input  [19:0] io_rxc_mem_0_c, 
  input  [19:0] io_rxc_mem_0_d, 
  input  [19:0] io_rxc_mem_0_e, 
  output        io_rxc_ridx, 
  input         io_rxc_widx, 
  output        io_rxc_safe_ridx_valid, 
  input         io_rxc_safe_widx_valid, 
  input         io_rxc_safe_source_reset_n, 
  output        io_rxc_safe_sink_reset_n, 
  input  [19:0] io_txc_mem_0_a, 
  input  [19:0] io_txc_mem_0_b, 
  input  [19:0] io_txc_mem_0_c, 
  input  [19:0] io_txc_mem_0_d, 
  input  [19:0] io_txc_mem_0_e, 
  output        io_txc_ridx, 
  input         io_txc_widx, 
  output        io_txc_safe_ridx_valid, 
  input         io_txc_safe_widx_valid, 
  input         io_txc_safe_source_reset_n, 
  output        io_txc_safe_sink_reset_n 
);
  wire  AsyncQueueSink_clock; 
  wire  AsyncQueueSink_reset; 
  wire  AsyncQueueSink_io_deq_ready; 
  wire  AsyncQueueSink_io_deq_valid; 
  wire [19:0] AsyncQueueSink_io_deq_bits_a; 
  wire [19:0] AsyncQueueSink_io_deq_bits_b; 
  wire [19:0] AsyncQueueSink_io_deq_bits_c; 
  wire [19:0] AsyncQueueSink_io_deq_bits_d; 
  wire [19:0] AsyncQueueSink_io_deq_bits_e; 
  wire [19:0] AsyncQueueSink_io_async_mem_0_a; 
  wire [19:0] AsyncQueueSink_io_async_mem_0_b; 
  wire [19:0] AsyncQueueSink_io_async_mem_0_c; 
  wire [19:0] AsyncQueueSink_io_async_mem_0_d; 
  wire [19:0] AsyncQueueSink_io_async_mem_0_e; 
  wire  AsyncQueueSink_io_async_ridx; 
  wire  AsyncQueueSink_io_async_widx; 
  wire  AsyncQueueSink_io_async_safe_ridx_valid; 
  wire  AsyncQueueSink_io_async_safe_widx_valid; 
  wire  AsyncQueueSink_io_async_safe_source_reset_n; 
  wire  AsyncQueueSink_io_async_safe_sink_reset_n; 
  wire  AsyncQueueSink_1_clock; 
  wire  AsyncQueueSink_1_reset; 
  wire  AsyncQueueSink_1_io_deq_ready; 
  wire  AsyncQueueSink_1_io_deq_valid; 
  wire [19:0] AsyncQueueSink_1_io_deq_bits_a; 
  wire [19:0] AsyncQueueSink_1_io_deq_bits_b; 
  wire [19:0] AsyncQueueSink_1_io_deq_bits_c; 
  wire [19:0] AsyncQueueSink_1_io_deq_bits_d; 
  wire [19:0] AsyncQueueSink_1_io_deq_bits_e; 
  wire [19:0] AsyncQueueSink_1_io_async_mem_0_a; 
  wire [19:0] AsyncQueueSink_1_io_async_mem_0_b; 
  wire [19:0] AsyncQueueSink_1_io_async_mem_0_c; 
  wire [19:0] AsyncQueueSink_1_io_async_mem_0_d; 
  wire [19:0] AsyncQueueSink_1_io_async_mem_0_e; 
  wire  AsyncQueueSink_1_io_async_ridx; 
  wire  AsyncQueueSink_1_io_async_widx; 
  wire  AsyncQueueSink_1_io_async_safe_ridx_valid; 
  wire  AsyncQueueSink_1_io_async_safe_widx_valid; 
  wire  AsyncQueueSink_1_io_async_safe_source_reset_n; 
  wire  AsyncQueueSink_1_io_async_safe_sink_reset_n; 
  wire  ShiftQueue_clock; 
  wire  ShiftQueue_reset; 
  wire  ShiftQueue_io_enq_ready; 
  wire  ShiftQueue_io_enq_valid; 
  wire [31:0] ShiftQueue_io_enq_bits_data; 
  wire  ShiftQueue_io_enq_bits_last; 
  wire [12:0] ShiftQueue_io_enq_bits_beats; 
  wire  ShiftQueue_io_deq_ready; 
  wire  ShiftQueue_io_deq_valid; 
  wire [31:0] ShiftQueue_io_deq_bits_data; 
  wire  ShiftQueue_io_deq_bits_last; 
  wire [12:0] ShiftQueue_io_deq_bits_beats; 
  wire  ShiftQueue_1_clock; 
  wire  ShiftQueue_1_reset; 
  wire  ShiftQueue_1_io_enq_ready; 
  wire  ShiftQueue_1_io_enq_valid; 
  wire [31:0] ShiftQueue_1_io_enq_bits_data; 
  wire  ShiftQueue_1_io_enq_bits_last; 
  wire [12:0] ShiftQueue_1_io_enq_bits_beats; 
  wire  ShiftQueue_1_io_deq_ready; 
  wire  ShiftQueue_1_io_deq_valid; 
  wire [31:0] ShiftQueue_1_io_deq_bits_data; 
  wire  ShiftQueue_1_io_deq_bits_last; 
  wire [12:0] ShiftQueue_1_io_deq_bits_beats; 
  wire  ShiftQueue_2_clock; 
  wire  ShiftQueue_2_reset; 
  wire  ShiftQueue_2_io_enq_ready; 
  wire  ShiftQueue_2_io_enq_valid; 
  wire [31:0] ShiftQueue_2_io_enq_bits_data; 
  wire  ShiftQueue_2_io_enq_bits_last; 
  wire [12:0] ShiftQueue_2_io_enq_bits_beats; 
  wire  ShiftQueue_2_io_deq_ready; 
  wire  ShiftQueue_2_io_deq_valid; 
  wire [31:0] ShiftQueue_2_io_deq_bits_data; 
  wire  ShiftQueue_2_io_deq_bits_last; 
  wire [12:0] ShiftQueue_2_io_deq_bits_beats; 
  wire  ShiftQueue_3_clock; 
  wire  ShiftQueue_3_reset; 
  wire  ShiftQueue_3_io_enq_ready; 
  wire  ShiftQueue_3_io_enq_valid; 
  wire [31:0] ShiftQueue_3_io_enq_bits_data; 
  wire  ShiftQueue_3_io_enq_bits_last; 
  wire [12:0] ShiftQueue_3_io_enq_bits_beats; 
  wire  ShiftQueue_3_io_deq_ready; 
  wire  ShiftQueue_3_io_deq_valid; 
  wire [31:0] ShiftQueue_3_io_deq_bits_data; 
  wire  ShiftQueue_3_io_deq_bits_last; 
  wire [12:0] ShiftQueue_3_io_deq_bits_beats; 
  wire  ShiftQueue_4_clock; 
  wire  ShiftQueue_4_reset; 
  wire  ShiftQueue_4_io_enq_ready; 
  wire  ShiftQueue_4_io_enq_valid; 
  wire [31:0] ShiftQueue_4_io_enq_bits_data; 
  wire  ShiftQueue_4_io_enq_bits_last; 
  wire [12:0] ShiftQueue_4_io_enq_bits_beats; 
  wire  ShiftQueue_4_io_deq_ready; 
  wire  ShiftQueue_4_io_deq_valid; 
  wire [31:0] ShiftQueue_4_io_deq_bits_data; 
  wire  ShiftQueue_4_io_deq_bits_last; 
  wire [12:0] ShiftQueue_4_io_deq_bits_beats; 
  wire  ShiftQueue_5_clock; 
  wire  ShiftQueue_5_reset; 
  wire  ShiftQueue_5_io_enq_ready; 
  wire  ShiftQueue_5_io_enq_valid; 
  wire [31:0] ShiftQueue_5_io_enq_bits_data; 
  wire  ShiftQueue_5_io_enq_bits_last; 
  wire [12:0] ShiftQueue_5_io_enq_bits_beats; 
  wire  ShiftQueue_5_io_deq_ready; 
  wire  ShiftQueue_5_io_deq_valid; 
  wire [31:0] ShiftQueue_5_io_deq_bits_data; 
  wire  ShiftQueue_5_io_deq_bits_last; 
  wire [12:0] ShiftQueue_5_io_deq_bits_beats; 
  wire  ShiftQueue_6_clock; 
  wire  ShiftQueue_6_reset; 
  wire  ShiftQueue_6_io_enq_ready; 
  wire  ShiftQueue_6_io_enq_valid; 
  wire [31:0] ShiftQueue_6_io_enq_bits_data; 
  wire  ShiftQueue_6_io_enq_bits_last; 
  wire [12:0] ShiftQueue_6_io_enq_bits_beats; 
  wire  ShiftQueue_6_io_deq_ready; 
  wire  ShiftQueue_6_io_deq_valid; 
  wire [31:0] ShiftQueue_6_io_deq_bits_data; 
  wire  ShiftQueue_6_io_deq_bits_last; 
  wire [12:0] ShiftQueue_6_io_deq_bits_beats; 
  wire  ShiftQueue_7_clock; 
  wire  ShiftQueue_7_reset; 
  wire  ShiftQueue_7_io_enq_ready; 
  wire  ShiftQueue_7_io_enq_valid; 
  wire [31:0] ShiftQueue_7_io_enq_bits_data; 
  wire  ShiftQueue_7_io_enq_bits_last; 
  wire [12:0] ShiftQueue_7_io_enq_bits_beats; 
  wire  ShiftQueue_7_io_deq_ready; 
  wire  ShiftQueue_7_io_deq_valid; 
  wire [31:0] ShiftQueue_7_io_deq_bits_data; 
  wire  ShiftQueue_7_io_deq_bits_last; 
  wire [12:0] ShiftQueue_7_io_deq_bits_beats; 
  wire  ShiftQueue_8_clock; 
  wire  ShiftQueue_8_reset; 
  wire  ShiftQueue_8_io_enq_ready; 
  wire  ShiftQueue_8_io_enq_valid; 
  wire [31:0] ShiftQueue_8_io_enq_bits_data; 
  wire  ShiftQueue_8_io_enq_bits_last; 
  wire [12:0] ShiftQueue_8_io_enq_bits_beats; 
  wire  ShiftQueue_8_io_deq_ready; 
  wire  ShiftQueue_8_io_deq_valid; 
  wire [31:0] ShiftQueue_8_io_deq_bits_data; 
  wire  ShiftQueue_8_io_deq_bits_last; 
  wire [12:0] ShiftQueue_8_io_deq_bits_beats; 
  wire  ShiftQueue_9_clock; 
  wire  ShiftQueue_9_reset; 
  wire  ShiftQueue_9_io_enq_ready; 
  wire  ShiftQueue_9_io_enq_valid; 
  wire [31:0] ShiftQueue_9_io_enq_bits_data; 
  wire  ShiftQueue_9_io_enq_bits_last; 
  wire [12:0] ShiftQueue_9_io_enq_bits_beats; 
  wire  ShiftQueue_9_io_deq_ready; 
  wire  ShiftQueue_9_io_deq_valid; 
  wire [31:0] ShiftQueue_9_io_deq_bits_data; 
  wire  ShiftQueue_9_io_deq_bits_last; 
  wire [12:0] ShiftQueue_9_io_deq_bits_beats; 
  wire  rxQ_clock; 
  wire  rxQ_reset; 
  wire  rxQ_io_enq_ready; 
  wire  rxQ_io_enq_valid; 
  wire [31:0] rxQ_io_enq_bits_data; 
  wire  rxQ_io_enq_bits_last; 
  wire [12:0] rxQ_io_enq_bits_beats; 
  wire  rxQ_io_deq_ready; 
  wire  rxQ_io_deq_valid; 
  wire [31:0] rxQ_io_deq_bits_data; 
  wire  rxQ_io_deq_bits_last; 
  wire [12:0] rxQ_io_deq_bits_beats; 
  wire  AsyncResetReg_d; 
  wire  AsyncResetReg_q; 
  wire  AsyncResetReg_en; 
  wire  AsyncResetReg_clk; 
  wire  AsyncResetReg_rst; 
  reg [19:0] rx_a; 
  reg [31:0] _RAND_0;
  reg [19:0] rx_b; 
  reg [31:0] _RAND_1;
  reg [19:0] rx_c; 
  reg [31:0] _RAND_2;
  reg [19:0] rx_d; 
  reg [31:0] _RAND_3;
  reg [19:0] rx_e; 
  reg [31:0] _RAND_4;
  reg [19:0] tx_a; 
  reg [31:0] _RAND_5;
  reg [19:0] tx_b; 
  reg [31:0] _RAND_6;
  reg [19:0] tx_c; 
  reg [31:0] _RAND_7;
  reg [19:0] tx_d; 
  reg [31:0] _RAND_8;
  reg [19:0] tx_e; 
  reg [31:0] _RAND_9;
  wire  _T_2; 
  reg  _T_3; 
  reg [31:0] _RAND_10;
  wire [19:0] _GEN_10; 
  wire [20:0] _T_4; 
  wire [20:0] _T_5; 
  wire  _T_6; 
  wire [20:0] _T_7; 
  wire  _T_8; 
  wire  _T_9; 
  wire  _T_11; 
  wire [20:0] _T_12; 
  wire  _T_13; 
  wire [19:0] _T_14; 
  wire [20:0] _GEN_11; 
  wire [20:0] _T_16; 
  wire  _T_19; 
  reg  _T_20; 
  reg [31:0] _RAND_11;
  wire [19:0] _GEN_12; 
  wire [20:0] _T_21; 
  wire [20:0] _T_22; 
  wire  _T_23; 
  wire [20:0] _T_24; 
  wire  _T_25; 
  wire  _T_26; 
  wire  _T_28; 
  wire [20:0] _T_29; 
  wire [19:0] _T_31; 
  wire [20:0] _GEN_13; 
  wire [20:0] _T_33; 
  wire  _T_36; 
  reg  _T_37; 
  reg [31:0] _RAND_12;
  wire [19:0] _GEN_14; 
  wire [20:0] _T_38; 
  wire [20:0] _T_39; 
  wire  _T_40; 
  wire [20:0] _T_41; 
  wire  _T_42; 
  wire  _T_43; 
  wire  _T_45; 
  wire [20:0] _T_46; 
  wire [19:0] _T_48; 
  wire [20:0] _GEN_15; 
  wire [20:0] _T_50; 
  wire  _T_53; 
  reg  _T_54; 
  reg [31:0] _RAND_13;
  wire [19:0] _GEN_16; 
  wire [20:0] _T_55; 
  wire [20:0] _T_56; 
  wire  _T_57; 
  wire [20:0] _T_58; 
  wire  _T_59; 
  wire  _T_60; 
  wire  _T_62; 
  wire [20:0] _T_63; 
  wire [19:0] _T_65; 
  wire [20:0] _GEN_17; 
  wire [20:0] _T_67; 
  wire  _T_70; 
  reg  _T_71; 
  reg [31:0] _RAND_14;
  wire [19:0] _GEN_18; 
  wire [20:0] _T_72; 
  wire [20:0] _T_73; 
  wire  _T_74; 
  wire [20:0] _T_75; 
  wire  _T_76; 
  wire  _T_77; 
  wire  _T_79; 
  wire [20:0] _T_80; 
  wire [19:0] _T_82; 
  wire [20:0] _GEN_19; 
  wire [20:0] _T_84; 
  wire [18:0] _T_87; 
  wire [19:0] _GEN_20; 
  wire [19:0] _T_88; 
  wire [17:0] _T_89; 
  wire [19:0] _GEN_21; 
  wire [19:0] _T_90; 
  wire [15:0] _T_91; 
  wire [19:0] _GEN_22; 
  wire [19:0] _T_92; 
  wire [11:0] _T_93; 
  wire [19:0] _GEN_23; 
  wire [19:0] _T_94; 
  wire [3:0] _T_95; 
  wire [19:0] _GEN_24; 
  wire [19:0] _T_96; 
  wire [18:0] _T_98; 
  wire [19:0] _T_99; 
  wire [19:0] _GEN_25; 
  wire [19:0] _T_100; 
  wire [19:0] _T_101; 
  wire [20:0] _T_102; 
  wire [4:0] _T_103; 
  wire [15:0] _T_104; 
  wire  _T_105; 
  wire [15:0] _GEN_26; 
  wire [15:0] _T_106; 
  wire [7:0] _T_107; 
  wire [7:0] _T_108; 
  wire  _T_109; 
  wire [7:0] _T_110; 
  wire [3:0] _T_111; 
  wire [3:0] _T_112; 
  wire  _T_113; 
  wire [3:0] _T_114; 
  wire [1:0] _T_115; 
  wire [1:0] _T_116; 
  wire  _T_117; 
  wire [1:0] _T_118; 
  wire  _T_119; 
  wire [19:0] rxLeft_a; 
  wire [18:0] _T_127; 
  wire [19:0] _GEN_28; 
  wire [19:0] _T_128; 
  wire [17:0] _T_129; 
  wire [19:0] _GEN_29; 
  wire [19:0] _T_130; 
  wire [15:0] _T_131; 
  wire [19:0] _GEN_30; 
  wire [19:0] _T_132; 
  wire [11:0] _T_133; 
  wire [19:0] _GEN_31; 
  wire [19:0] _T_134; 
  wire [3:0] _T_135; 
  wire [19:0] _GEN_32; 
  wire [19:0] _T_136; 
  wire [18:0] _T_138; 
  wire [19:0] _T_139; 
  wire [19:0] _GEN_33; 
  wire [19:0] _T_140; 
  wire [19:0] _T_141; 
  wire [20:0] _T_142; 
  wire [4:0] _T_143; 
  wire [15:0] _T_144; 
  wire  _T_145; 
  wire [15:0] _GEN_34; 
  wire [15:0] _T_146; 
  wire [7:0] _T_147; 
  wire [7:0] _T_148; 
  wire  _T_149; 
  wire [7:0] _T_150; 
  wire [3:0] _T_151; 
  wire [3:0] _T_152; 
  wire  _T_153; 
  wire [3:0] _T_154; 
  wire [1:0] _T_155; 
  wire [1:0] _T_156; 
  wire  _T_157; 
  wire [1:0] _T_158; 
  wire  _T_159; 
  wire [19:0] rxLeft_b; 
  wire [18:0] _T_167; 
  wire [19:0] _GEN_36; 
  wire [19:0] _T_168; 
  wire [17:0] _T_169; 
  wire [19:0] _GEN_37; 
  wire [19:0] _T_170; 
  wire [15:0] _T_171; 
  wire [19:0] _GEN_38; 
  wire [19:0] _T_172; 
  wire [11:0] _T_173; 
  wire [19:0] _GEN_39; 
  wire [19:0] _T_174; 
  wire [3:0] _T_175; 
  wire [19:0] _GEN_40; 
  wire [19:0] _T_176; 
  wire [18:0] _T_178; 
  wire [19:0] _T_179; 
  wire [19:0] _GEN_41; 
  wire [19:0] _T_180; 
  wire [19:0] _T_181; 
  wire [20:0] _T_182; 
  wire [4:0] _T_183; 
  wire [15:0] _T_184; 
  wire  _T_185; 
  wire [15:0] _GEN_42; 
  wire [15:0] _T_186; 
  wire [7:0] _T_187; 
  wire [7:0] _T_188; 
  wire  _T_189; 
  wire [7:0] _T_190; 
  wire [3:0] _T_191; 
  wire [3:0] _T_192; 
  wire  _T_193; 
  wire [3:0] _T_194; 
  wire [1:0] _T_195; 
  wire [1:0] _T_196; 
  wire  _T_197; 
  wire [1:0] _T_198; 
  wire  _T_199; 
  wire [19:0] rxLeft_c; 
  wire [18:0] _T_207; 
  wire [19:0] _GEN_44; 
  wire [19:0] _T_208; 
  wire [17:0] _T_209; 
  wire [19:0] _GEN_45; 
  wire [19:0] _T_210; 
  wire [15:0] _T_211; 
  wire [19:0] _GEN_46; 
  wire [19:0] _T_212; 
  wire [11:0] _T_213; 
  wire [19:0] _GEN_47; 
  wire [19:0] _T_214; 
  wire [3:0] _T_215; 
  wire [19:0] _GEN_48; 
  wire [19:0] _T_216; 
  wire [18:0] _T_218; 
  wire [19:0] _T_219; 
  wire [19:0] _GEN_49; 
  wire [19:0] _T_220; 
  wire [19:0] _T_221; 
  wire [20:0] _T_222; 
  wire [4:0] _T_223; 
  wire [15:0] _T_224; 
  wire  _T_225; 
  wire [15:0] _GEN_50; 
  wire [15:0] _T_226; 
  wire [7:0] _T_227; 
  wire [7:0] _T_228; 
  wire  _T_229; 
  wire [7:0] _T_230; 
  wire [3:0] _T_231; 
  wire [3:0] _T_232; 
  wire  _T_233; 
  wire [3:0] _T_234; 
  wire [1:0] _T_235; 
  wire [1:0] _T_236; 
  wire  _T_237; 
  wire [1:0] _T_238; 
  wire  _T_239; 
  wire [19:0] rxLeft_d; 
  wire [18:0] _T_247; 
  wire [19:0] _GEN_52; 
  wire [19:0] _T_248; 
  wire [17:0] _T_249; 
  wire [19:0] _GEN_53; 
  wire [19:0] _T_250; 
  wire [15:0] _T_251; 
  wire [19:0] _GEN_54; 
  wire [19:0] _T_252; 
  wire [11:0] _T_253; 
  wire [19:0] _GEN_55; 
  wire [19:0] _T_254; 
  wire [3:0] _T_255; 
  wire [19:0] _GEN_56; 
  wire [19:0] _T_256; 
  wire [18:0] _T_258; 
  wire [19:0] _T_259; 
  wire [19:0] _GEN_57; 
  wire [19:0] _T_260; 
  wire [19:0] _T_261; 
  wire [20:0] _T_262; 
  wire [4:0] _T_263; 
  wire [15:0] _T_264; 
  wire  _T_265; 
  wire [15:0] _GEN_58; 
  wire [15:0] _T_266; 
  wire [7:0] _T_267; 
  wire [7:0] _T_268; 
  wire  _T_269; 
  wire [7:0] _T_270; 
  wire [3:0] _T_271; 
  wire [3:0] _T_272; 
  wire  _T_273; 
  wire [3:0] _T_274; 
  wire [1:0] _T_275; 
  wire [1:0] _T_276; 
  wire  _T_277; 
  wire [1:0] _T_278; 
  wire  _T_279; 
  wire [19:0] rxLeft_e; 
  wire [11:0] _T_288; 
  wire [9:0] _T_289; 
  wire [9:0] _T_290; 
  wire [19:0] _T_291; 
  wire  _T_292; 
  wire [19:0] _T_293_a; 
  wire [19:0] _T_293_b; 
  wire [19:0] _T_293_c; 
  wire [19:0] _T_293_d; 
  wire [19:0] _T_293_e; 
  wire  _T_294; 
  wire [19:0] _T_296_a; 
  wire [19:0] _T_296_b; 
  wire [19:0] _T_296_c; 
  wire [19:0] _T_296_d; 
  wire [19:0] _T_296_e; 
  wire [20:0] _T_298; 
  wire  _T_299; 
  wire [20:0] _T_302; 
  wire [20:0] _T_303; 
  wire  _T_304; 
  wire [20:0] _T_307; 
  wire [20:0] _T_308; 
  wire  _T_309; 
  wire [20:0] _T_312; 
  wire [20:0] _T_313; 
  wire  _T_314; 
  wire [20:0] _T_317; 
  wire [20:0] _T_318; 
  wire  _T_319; 
  wire [20:0] _T_322; 
  wire  _T_336; 
  wire  _T_337; 
  wire  _T_338; 
  wire  _T_339; 
  wire  _T_340; 
  reg [4:0] xmit; 
  reg [31:0] _RAND_15;
  wire  forceXmit; 
  wire  allowReturn; 
  wire  f_valid; 
  wire [5:0] requests; 
  wire  f_bits_last; 
  wire [5:0] lasts; 
  wire  _T_331; 
  wire [4:0] _T_333; 
  reg  first; 
  reg [31:0] _RAND_16;
  reg [5:0] _T_349; 
  reg [31:0] _RAND_17;
  wire [5:0] _T_350; 
  wire [5:0] _T_351; 
  wire [11:0] _T_352; 
  wire [10:0] _T_353; 
  wire [11:0] _GEN_60; 
  wire [11:0] _T_354; 
  wire [9:0] _T_355; 
  wire [11:0] _GEN_61; 
  wire [11:0] _T_356; 
  wire [7:0] _T_357; 
  wire [11:0] _GEN_62; 
  wire [11:0] _T_358; 
  wire [10:0] _T_360; 
  wire [11:0] _T_361; 
  wire [11:0] _GEN_63; 
  wire [11:0] _T_362; 
  wire [5:0] _T_363; 
  wire [5:0] _T_364; 
  wire [5:0] _T_365; 
  wire [5:0] readys; 
  reg [5:0] state; 
  reg [31:0] _RAND_18;
  wire [5:0] allowed; 
  wire  f_ready; 
  wire  _T_334; 
  wire  _T_344; 
  wire  _T_346; 
  wire  _T_347; 
  wire  _T_367; 
  wire  _T_368; 
  wire [5:0] _T_369; 
  wire [6:0] _T_370; 
  wire [5:0] _T_371; 
  wire [5:0] _T_372; 
  wire [7:0] _T_373; 
  wire [5:0] _T_374; 
  wire [5:0] _T_375; 
  wire [9:0] _T_376; 
  wire [5:0] _T_377; 
  wire [5:0] _T_378; 
  wire [5:0] grant; 
  wire [5:0] _T_386; 
  wire  _T_387; 
  wire  send; 
  wire [5:0] _T_388; 
  wire  _T_389; 
  wire  _T_390; 
  wire  _T_392; 
  wire  _T_393; 
  wire [5:0] _T_394; 
  wire  _T_395; 
  reg  _T_397; 
  reg [31:0] _RAND_19;
  reg  _T_398; 
  reg [31:0] _RAND_20;
  reg [5:0] _T_399; 
  reg [31:0] _RAND_21;
  reg [31:0] _T_401_0; 
  reg [31:0] _RAND_22;
  reg [31:0] _T_401_1; 
  reg [31:0] _RAND_23;
  reg [31:0] _T_401_2; 
  reg [31:0] _RAND_24;
  reg [31:0] _T_401_3; 
  reg [31:0] _RAND_25;
  reg [31:0] _T_401_4; 
  reg [31:0] _RAND_26;
  reg [31:0] _T_401_5; 
  reg [31:0] _RAND_27;
  wire  _T_402; 
  wire  _T_403; 
  wire  _T_404; 
  wire  _T_405; 
  wire  _T_406; 
  wire  _T_407; 
  wire [31:0] _T_408; 
  wire [31:0] _T_409; 
  wire [31:0] _T_410; 
  wire [31:0] _T_411; 
  wire [31:0] _T_412; 
  wire [31:0] _T_413; 
  wire [31:0] _T_414; 
  wire [31:0] _T_415; 
  wire [31:0] _T_416; 
  wire [31:0] _T_417; 
  reg [31:0] _T_420; 
  reg [31:0] _RAND_28;
  wire [19:0] _T_297_a; 
  wire [19:0] _T_297_b; 
  wire [19:0] _T_297_c; 
  wire [19:0] _T_297_d; 
  wire [19:0] _T_297_e; 
  dual_AsyncQueueSink_5 dual_AsyncQueueSink ( 
    .clock(AsyncQueueSink_clock),
    .reset(AsyncQueueSink_reset),
    .io_deq_ready(AsyncQueueSink_io_deq_ready),
    .io_deq_valid(AsyncQueueSink_io_deq_valid),
    .io_deq_bits_a(AsyncQueueSink_io_deq_bits_a),
    .io_deq_bits_b(AsyncQueueSink_io_deq_bits_b),
    .io_deq_bits_c(AsyncQueueSink_io_deq_bits_c),
    .io_deq_bits_d(AsyncQueueSink_io_deq_bits_d),
    .io_deq_bits_e(AsyncQueueSink_io_deq_bits_e),
    .io_async_mem_0_a(AsyncQueueSink_io_async_mem_0_a),
    .io_async_mem_0_b(AsyncQueueSink_io_async_mem_0_b),
    .io_async_mem_0_c(AsyncQueueSink_io_async_mem_0_c),
    .io_async_mem_0_d(AsyncQueueSink_io_async_mem_0_d),
    .io_async_mem_0_e(AsyncQueueSink_io_async_mem_0_e),
    .io_async_ridx(AsyncQueueSink_io_async_ridx),
    .io_async_widx(AsyncQueueSink_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSink_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSink_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSink_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSink_io_async_safe_sink_reset_n)
  );
  dual_AsyncQueueSink_5 AsyncQueueSink_1 ( 
    .clock(AsyncQueueSink_1_clock),
    .reset(AsyncQueueSink_1_reset),
    .io_deq_ready(AsyncQueueSink_1_io_deq_ready),
    .io_deq_valid(AsyncQueueSink_1_io_deq_valid),
    .io_deq_bits_a(AsyncQueueSink_1_io_deq_bits_a),
    .io_deq_bits_b(AsyncQueueSink_1_io_deq_bits_b),
    .io_deq_bits_c(AsyncQueueSink_1_io_deq_bits_c),
    .io_deq_bits_d(AsyncQueueSink_1_io_deq_bits_d),
    .io_deq_bits_e(AsyncQueueSink_1_io_deq_bits_e),
    .io_async_mem_0_a(AsyncQueueSink_1_io_async_mem_0_a),
    .io_async_mem_0_b(AsyncQueueSink_1_io_async_mem_0_b),
    .io_async_mem_0_c(AsyncQueueSink_1_io_async_mem_0_c),
    .io_async_mem_0_d(AsyncQueueSink_1_io_async_mem_0_d),
    .io_async_mem_0_e(AsyncQueueSink_1_io_async_mem_0_e),
    .io_async_ridx(AsyncQueueSink_1_io_async_ridx),
    .io_async_widx(AsyncQueueSink_1_io_async_widx),
    .io_async_safe_ridx_valid(AsyncQueueSink_1_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(AsyncQueueSink_1_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(AsyncQueueSink_1_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(AsyncQueueSink_1_io_async_safe_sink_reset_n)
  );
  dual_ShiftQueue ShiftQueue ( 
    .clock(ShiftQueue_clock),
    .reset(ShiftQueue_reset),
    .io_enq_ready(ShiftQueue_io_enq_ready),
    .io_enq_valid(ShiftQueue_io_enq_valid),
    .io_enq_bits_data(ShiftQueue_io_enq_bits_data),
    .io_enq_bits_last(ShiftQueue_io_enq_bits_last),
    .io_enq_bits_beats(ShiftQueue_io_enq_bits_beats),
    .io_deq_ready(ShiftQueue_io_deq_ready),
    .io_deq_valid(ShiftQueue_io_deq_valid),
    .io_deq_bits_data(ShiftQueue_io_deq_bits_data),
    .io_deq_bits_last(ShiftQueue_io_deq_bits_last),
    .io_deq_bits_beats(ShiftQueue_io_deq_bits_beats)
  );
  dual_ShiftQueue ShiftQueue_1 ( 
    .clock(ShiftQueue_1_clock),
    .reset(ShiftQueue_1_reset),
    .io_enq_ready(ShiftQueue_1_io_enq_ready),
    .io_enq_valid(ShiftQueue_1_io_enq_valid),
    .io_enq_bits_data(ShiftQueue_1_io_enq_bits_data),
    .io_enq_bits_last(ShiftQueue_1_io_enq_bits_last),
    .io_enq_bits_beats(ShiftQueue_1_io_enq_bits_beats),
    .io_deq_ready(ShiftQueue_1_io_deq_ready),
    .io_deq_valid(ShiftQueue_1_io_deq_valid),
    .io_deq_bits_data(ShiftQueue_1_io_deq_bits_data),
    .io_deq_bits_last(ShiftQueue_1_io_deq_bits_last),
    .io_deq_bits_beats(ShiftQueue_1_io_deq_bits_beats)
  );
  dual_ShiftQueue ShiftQueue_2 ( 
    .clock(ShiftQueue_2_clock),
    .reset(ShiftQueue_2_reset),
    .io_enq_ready(ShiftQueue_2_io_enq_ready),
    .io_enq_valid(ShiftQueue_2_io_enq_valid),
    .io_enq_bits_data(ShiftQueue_2_io_enq_bits_data),
    .io_enq_bits_last(ShiftQueue_2_io_enq_bits_last),
    .io_enq_bits_beats(ShiftQueue_2_io_enq_bits_beats),
    .io_deq_ready(ShiftQueue_2_io_deq_ready),
    .io_deq_valid(ShiftQueue_2_io_deq_valid),
    .io_deq_bits_data(ShiftQueue_2_io_deq_bits_data),
    .io_deq_bits_last(ShiftQueue_2_io_deq_bits_last),
    .io_deq_bits_beats(ShiftQueue_2_io_deq_bits_beats)
  );
  dual_ShiftQueue ShiftQueue_3 ( 
    .clock(ShiftQueue_3_clock),
    .reset(ShiftQueue_3_reset),
    .io_enq_ready(ShiftQueue_3_io_enq_ready),
    .io_enq_valid(ShiftQueue_3_io_enq_valid),
    .io_enq_bits_data(ShiftQueue_3_io_enq_bits_data),
    .io_enq_bits_last(ShiftQueue_3_io_enq_bits_last),
    .io_enq_bits_beats(ShiftQueue_3_io_enq_bits_beats),
    .io_deq_ready(ShiftQueue_3_io_deq_ready),
    .io_deq_valid(ShiftQueue_3_io_deq_valid),
    .io_deq_bits_data(ShiftQueue_3_io_deq_bits_data),
    .io_deq_bits_last(ShiftQueue_3_io_deq_bits_last),
    .io_deq_bits_beats(ShiftQueue_3_io_deq_bits_beats)
  );
  dual_ShiftQueue ShiftQueue_4 ( 
    .clock(ShiftQueue_4_clock),
    .reset(ShiftQueue_4_reset),
    .io_enq_ready(ShiftQueue_4_io_enq_ready),
    .io_enq_valid(ShiftQueue_4_io_enq_valid),
    .io_enq_bits_data(ShiftQueue_4_io_enq_bits_data),
    .io_enq_bits_last(ShiftQueue_4_io_enq_bits_last),
    .io_enq_bits_beats(ShiftQueue_4_io_enq_bits_beats),
    .io_deq_ready(ShiftQueue_4_io_deq_ready),
    .io_deq_valid(ShiftQueue_4_io_deq_valid),
    .io_deq_bits_data(ShiftQueue_4_io_deq_bits_data),
    .io_deq_bits_last(ShiftQueue_4_io_deq_bits_last),
    .io_deq_bits_beats(ShiftQueue_4_io_deq_bits_beats)
  );
  dual_ShiftQueue ShiftQueue_5 ( 
    .clock(ShiftQueue_5_clock),
    .reset(ShiftQueue_5_reset),
    .io_enq_ready(ShiftQueue_5_io_enq_ready),
    .io_enq_valid(ShiftQueue_5_io_enq_valid),
    .io_enq_bits_data(ShiftQueue_5_io_enq_bits_data),
    .io_enq_bits_last(ShiftQueue_5_io_enq_bits_last),
    .io_enq_bits_beats(ShiftQueue_5_io_enq_bits_beats),
    .io_deq_ready(ShiftQueue_5_io_deq_ready),
    .io_deq_valid(ShiftQueue_5_io_deq_valid),
    .io_deq_bits_data(ShiftQueue_5_io_deq_bits_data),
    .io_deq_bits_last(ShiftQueue_5_io_deq_bits_last),
    .io_deq_bits_beats(ShiftQueue_5_io_deq_bits_beats)
  );
  dual_ShiftQueue ShiftQueue_6 ( 
    .clock(ShiftQueue_6_clock),
    .reset(ShiftQueue_6_reset),
    .io_enq_ready(ShiftQueue_6_io_enq_ready),
    .io_enq_valid(ShiftQueue_6_io_enq_valid),
    .io_enq_bits_data(ShiftQueue_6_io_enq_bits_data),
    .io_enq_bits_last(ShiftQueue_6_io_enq_bits_last),
    .io_enq_bits_beats(ShiftQueue_6_io_enq_bits_beats),
    .io_deq_ready(ShiftQueue_6_io_deq_ready),
    .io_deq_valid(ShiftQueue_6_io_deq_valid),
    .io_deq_bits_data(ShiftQueue_6_io_deq_bits_data),
    .io_deq_bits_last(ShiftQueue_6_io_deq_bits_last),
    .io_deq_bits_beats(ShiftQueue_6_io_deq_bits_beats)
  );
  dual_ShiftQueue ShiftQueue_7 ( 
    .clock(ShiftQueue_7_clock),
    .reset(ShiftQueue_7_reset),
    .io_enq_ready(ShiftQueue_7_io_enq_ready),
    .io_enq_valid(ShiftQueue_7_io_enq_valid),
    .io_enq_bits_data(ShiftQueue_7_io_enq_bits_data),
    .io_enq_bits_last(ShiftQueue_7_io_enq_bits_last),
    .io_enq_bits_beats(ShiftQueue_7_io_enq_bits_beats),
    .io_deq_ready(ShiftQueue_7_io_deq_ready),
    .io_deq_valid(ShiftQueue_7_io_deq_valid),
    .io_deq_bits_data(ShiftQueue_7_io_deq_bits_data),
    .io_deq_bits_last(ShiftQueue_7_io_deq_bits_last),
    .io_deq_bits_beats(ShiftQueue_7_io_deq_bits_beats)
  );
  dual_ShiftQueue ShiftQueue_8 ( 
    .clock(ShiftQueue_8_clock),
    .reset(ShiftQueue_8_reset),
    .io_enq_ready(ShiftQueue_8_io_enq_ready),
    .io_enq_valid(ShiftQueue_8_io_enq_valid),
    .io_enq_bits_data(ShiftQueue_8_io_enq_bits_data),
    .io_enq_bits_last(ShiftQueue_8_io_enq_bits_last),
    .io_enq_bits_beats(ShiftQueue_8_io_enq_bits_beats),
    .io_deq_ready(ShiftQueue_8_io_deq_ready),
    .io_deq_valid(ShiftQueue_8_io_deq_valid),
    .io_deq_bits_data(ShiftQueue_8_io_deq_bits_data),
    .io_deq_bits_last(ShiftQueue_8_io_deq_bits_last),
    .io_deq_bits_beats(ShiftQueue_8_io_deq_bits_beats)
  );
  dual_ShiftQueue ShiftQueue_9 ( 
    .clock(ShiftQueue_9_clock),
    .reset(ShiftQueue_9_reset),
    .io_enq_ready(ShiftQueue_9_io_enq_ready),
    .io_enq_valid(ShiftQueue_9_io_enq_valid),
    .io_enq_bits_data(ShiftQueue_9_io_enq_bits_data),
    .io_enq_bits_last(ShiftQueue_9_io_enq_bits_last),
    .io_enq_bits_beats(ShiftQueue_9_io_enq_bits_beats),
    .io_deq_ready(ShiftQueue_9_io_deq_ready),
    .io_deq_valid(ShiftQueue_9_io_deq_valid),
    .io_deq_bits_data(ShiftQueue_9_io_deq_bits_data),
    .io_deq_bits_last(ShiftQueue_9_io_deq_bits_last),
    .io_deq_bits_beats(ShiftQueue_9_io_deq_bits_beats)
  );
  dual_ShiftQueue rxQ ( 
    .clock(rxQ_clock),
    .reset(rxQ_reset),
    .io_enq_ready(rxQ_io_enq_ready),
    .io_enq_valid(rxQ_io_enq_valid),
    .io_enq_bits_data(rxQ_io_enq_bits_data),
    .io_enq_bits_last(rxQ_io_enq_bits_last),
    .io_enq_bits_beats(rxQ_io_enq_bits_beats),
    .io_deq_ready(rxQ_io_deq_ready),
    .io_deq_valid(rxQ_io_deq_valid),
    .io_deq_bits_data(rxQ_io_deq_bits_data),
    .io_deq_bits_last(rxQ_io_deq_bits_last),
    .io_deq_bits_beats(rxQ_io_deq_bits_beats)
  );
  dual_AsyncResetReg #(.RESET_VALUE(1)) AsyncResetReg ( 
    .d(AsyncResetReg_d),
    .q(AsyncResetReg_q),
    .en(AsyncResetReg_en),
    .clk(AsyncResetReg_clk),
    .rst(AsyncResetReg_rst)
  );
  assign _T_2 = ShiftQueue_io_deq_ready & ShiftQueue_io_deq_valid; 
  assign _GEN_10 = {{7'd0}, ShiftQueue_io_deq_bits_beats}; 
  assign _T_4 = tx_a - _GEN_10; 
  assign _T_5 = $unsigned(_T_4); 
  assign _T_6 = _T_3 == 1'h0; 
  assign _T_7 = $signed(_T_5); 
  assign _T_8 = $signed(_T_7) >= $signed(21'sh0); 
  assign _T_9 = _T_6 | _T_8; 
  assign _T_11 = _T_2 & _T_3; 
  assign _T_12 = _T_11 ? _T_5 : {{1'd0}, tx_a}; 
  assign _T_13 = AsyncQueueSink_1_io_deq_ready & AsyncQueueSink_1_io_deq_valid; 
  assign _T_14 = _T_13 ? AsyncQueueSink_1_io_deq_bits_a : 20'h0; 
  assign _GEN_11 = {{1'd0}, _T_14}; 
  assign _T_16 = _T_12 + _GEN_11; 
  assign _T_19 = ShiftQueue_1_io_deq_ready & ShiftQueue_1_io_deq_valid; 
  assign _GEN_12 = {{7'd0}, ShiftQueue_1_io_deq_bits_beats}; 
  assign _T_21 = tx_b - _GEN_12; 
  assign _T_22 = $unsigned(_T_21); 
  assign _T_23 = _T_20 == 1'h0; 
  assign _T_24 = $signed(_T_22); 
  assign _T_25 = $signed(_T_24) >= $signed(21'sh0); 
  assign _T_26 = _T_23 | _T_25; 
  assign _T_28 = _T_19 & _T_20; 
  assign _T_29 = _T_28 ? _T_22 : {{1'd0}, tx_b}; 
  assign _T_31 = _T_13 ? AsyncQueueSink_1_io_deq_bits_b : 20'h0; 
  assign _GEN_13 = {{1'd0}, _T_31}; 
  assign _T_33 = _T_29 + _GEN_13; 
  assign _T_36 = ShiftQueue_2_io_deq_ready & ShiftQueue_2_io_deq_valid; 
  assign _GEN_14 = {{7'd0}, ShiftQueue_2_io_deq_bits_beats}; 
  assign _T_38 = tx_c - _GEN_14; 
  assign _T_39 = $unsigned(_T_38); 
  assign _T_40 = _T_37 == 1'h0; 
  assign _T_41 = $signed(_T_39); 
  assign _T_42 = $signed(_T_41) >= $signed(21'sh0); 
  assign _T_43 = _T_40 | _T_42; 
  assign _T_45 = _T_36 & _T_37; 
  assign _T_46 = _T_45 ? _T_39 : {{1'd0}, tx_c}; 
  assign _T_48 = _T_13 ? AsyncQueueSink_1_io_deq_bits_c : 20'h0; 
  assign _GEN_15 = {{1'd0}, _T_48}; 
  assign _T_50 = _T_46 + _GEN_15; 
  assign _T_53 = ShiftQueue_3_io_deq_ready & ShiftQueue_3_io_deq_valid; 
  assign _GEN_16 = {{7'd0}, ShiftQueue_3_io_deq_bits_beats}; 
  assign _T_55 = tx_d - _GEN_16; 
  assign _T_56 = $unsigned(_T_55); 
  assign _T_57 = _T_54 == 1'h0; 
  assign _T_58 = $signed(_T_56); 
  assign _T_59 = $signed(_T_58) >= $signed(21'sh0); 
  assign _T_60 = _T_57 | _T_59; 
  assign _T_62 = _T_53 & _T_54; 
  assign _T_63 = _T_62 ? _T_56 : {{1'd0}, tx_d}; 
  assign _T_65 = _T_13 ? AsyncQueueSink_1_io_deq_bits_d : 20'h0; 
  assign _GEN_17 = {{1'd0}, _T_65}; 
  assign _T_67 = _T_63 + _GEN_17; 
  assign _T_70 = ShiftQueue_4_io_deq_ready & ShiftQueue_4_io_deq_valid; 
  assign _GEN_18 = {{7'd0}, ShiftQueue_4_io_deq_bits_beats}; 
  assign _T_72 = tx_e - _GEN_18; 
  assign _T_73 = $unsigned(_T_72); 
  assign _T_74 = _T_71 == 1'h0; 
  assign _T_75 = $signed(_T_73); 
  assign _T_76 = $signed(_T_75) >= $signed(21'sh0); 
  assign _T_77 = _T_74 | _T_76; 
  assign _T_79 = _T_70 & _T_71; 
  assign _T_80 = _T_79 ? _T_73 : {{1'd0}, tx_e}; 
  assign _T_82 = _T_13 ? AsyncQueueSink_1_io_deq_bits_e : 20'h0; 
  assign _GEN_19 = {{1'd0}, _T_82}; 
  assign _T_84 = _T_80 + _GEN_19; 
  assign _T_87 = rx_a[19:1]; 
  assign _GEN_20 = {{1'd0}, _T_87}; 
  assign _T_88 = rx_a | _GEN_20; 
  assign _T_89 = _T_88[19:2]; 
  assign _GEN_21 = {{2'd0}, _T_89}; 
  assign _T_90 = _T_88 | _GEN_21; 
  assign _T_91 = _T_90[19:4]; 
  assign _GEN_22 = {{4'd0}, _T_91}; 
  assign _T_92 = _T_90 | _GEN_22; 
  assign _T_93 = _T_92[19:8]; 
  assign _GEN_23 = {{8'd0}, _T_93}; 
  assign _T_94 = _T_92 | _GEN_23; 
  assign _T_95 = _T_94[19:16]; 
  assign _GEN_24 = {{16'd0}, _T_95}; 
  assign _T_96 = _T_94 | _GEN_24; 
  assign _T_98 = _T_96[19:1]; 
  assign _T_99 = ~ rx_a; 
  assign _GEN_25 = {{1'd0}, _T_98}; 
  assign _T_100 = _T_99 | _GEN_25; 
  assign _T_101 = ~ _T_100; 
  assign _T_102 = {_T_101, 1'h0}; 
  assign _T_103 = _T_102[20:16]; 
  assign _T_104 = _T_102[15:0]; 
  assign _T_105 = _T_103 != 5'h0; 
  assign _GEN_26 = {{11'd0}, _T_103}; 
  assign _T_106 = _GEN_26 | _T_104; 
  assign _T_107 = _T_106[15:8]; 
  assign _T_108 = _T_106[7:0]; 
  assign _T_109 = _T_107 != 8'h0; 
  assign _T_110 = _T_107 | _T_108; 
  assign _T_111 = _T_110[7:4]; 
  assign _T_112 = _T_110[3:0]; 
  assign _T_113 = _T_111 != 4'h0; 
  assign _T_114 = _T_111 | _T_112; 
  assign _T_115 = _T_114[3:2]; 
  assign _T_116 = _T_114[1:0]; 
  assign _T_117 = _T_115 != 2'h0; 
  assign _T_118 = _T_115 | _T_116; 
  assign _T_119 = _T_118[1]; 
  assign rxLeft_a = rx_a & _GEN_25; 
  assign _T_127 = rx_b[19:1]; 
  assign _GEN_28 = {{1'd0}, _T_127}; 
  assign _T_128 = rx_b | _GEN_28; 
  assign _T_129 = _T_128[19:2]; 
  assign _GEN_29 = {{2'd0}, _T_129}; 
  assign _T_130 = _T_128 | _GEN_29; 
  assign _T_131 = _T_130[19:4]; 
  assign _GEN_30 = {{4'd0}, _T_131}; 
  assign _T_132 = _T_130 | _GEN_30; 
  assign _T_133 = _T_132[19:8]; 
  assign _GEN_31 = {{8'd0}, _T_133}; 
  assign _T_134 = _T_132 | _GEN_31; 
  assign _T_135 = _T_134[19:16]; 
  assign _GEN_32 = {{16'd0}, _T_135}; 
  assign _T_136 = _T_134 | _GEN_32; 
  assign _T_138 = _T_136[19:1]; 
  assign _T_139 = ~ rx_b; 
  assign _GEN_33 = {{1'd0}, _T_138}; 
  assign _T_140 = _T_139 | _GEN_33; 
  assign _T_141 = ~ _T_140; 
  assign _T_142 = {_T_141, 1'h0}; 
  assign _T_143 = _T_142[20:16]; 
  assign _T_144 = _T_142[15:0]; 
  assign _T_145 = _T_143 != 5'h0; 
  assign _GEN_34 = {{11'd0}, _T_143}; 
  assign _T_146 = _GEN_34 | _T_144; 
  assign _T_147 = _T_146[15:8]; 
  assign _T_148 = _T_146[7:0]; 
  assign _T_149 = _T_147 != 8'h0; 
  assign _T_150 = _T_147 | _T_148; 
  assign _T_151 = _T_150[7:4]; 
  assign _T_152 = _T_150[3:0]; 
  assign _T_153 = _T_151 != 4'h0; 
  assign _T_154 = _T_151 | _T_152; 
  assign _T_155 = _T_154[3:2]; 
  assign _T_156 = _T_154[1:0]; 
  assign _T_157 = _T_155 != 2'h0; 
  assign _T_158 = _T_155 | _T_156; 
  assign _T_159 = _T_158[1]; 
  assign rxLeft_b = rx_b & _GEN_33; 
  assign _T_167 = rx_c[19:1]; 
  assign _GEN_36 = {{1'd0}, _T_167}; 
  assign _T_168 = rx_c | _GEN_36; 
  assign _T_169 = _T_168[19:2]; 
  assign _GEN_37 = {{2'd0}, _T_169}; 
  assign _T_170 = _T_168 | _GEN_37; 
  assign _T_171 = _T_170[19:4]; 
  assign _GEN_38 = {{4'd0}, _T_171}; 
  assign _T_172 = _T_170 | _GEN_38; 
  assign _T_173 = _T_172[19:8]; 
  assign _GEN_39 = {{8'd0}, _T_173}; 
  assign _T_174 = _T_172 | _GEN_39; 
  assign _T_175 = _T_174[19:16]; 
  assign _GEN_40 = {{16'd0}, _T_175}; 
  assign _T_176 = _T_174 | _GEN_40; 
  assign _T_178 = _T_176[19:1]; 
  assign _T_179 = ~ rx_c; 
  assign _GEN_41 = {{1'd0}, _T_178}; 
  assign _T_180 = _T_179 | _GEN_41; 
  assign _T_181 = ~ _T_180; 
  assign _T_182 = {_T_181, 1'h0}; 
  assign _T_183 = _T_182[20:16]; 
  assign _T_184 = _T_182[15:0]; 
  assign _T_185 = _T_183 != 5'h0; 
  assign _GEN_42 = {{11'd0}, _T_183}; 
  assign _T_186 = _GEN_42 | _T_184; 
  assign _T_187 = _T_186[15:8]; 
  assign _T_188 = _T_186[7:0]; 
  assign _T_189 = _T_187 != 8'h0; 
  assign _T_190 = _T_187 | _T_188; 
  assign _T_191 = _T_190[7:4]; 
  assign _T_192 = _T_190[3:0]; 
  assign _T_193 = _T_191 != 4'h0; 
  assign _T_194 = _T_191 | _T_192; 
  assign _T_195 = _T_194[3:2]; 
  assign _T_196 = _T_194[1:0]; 
  assign _T_197 = _T_195 != 2'h0; 
  assign _T_198 = _T_195 | _T_196; 
  assign _T_199 = _T_198[1]; 
  assign rxLeft_c = rx_c & _GEN_41; 
  assign _T_207 = rx_d[19:1]; 
  assign _GEN_44 = {{1'd0}, _T_207}; 
  assign _T_208 = rx_d | _GEN_44; 
  assign _T_209 = _T_208[19:2]; 
  assign _GEN_45 = {{2'd0}, _T_209}; 
  assign _T_210 = _T_208 | _GEN_45; 
  assign _T_211 = _T_210[19:4]; 
  assign _GEN_46 = {{4'd0}, _T_211}; 
  assign _T_212 = _T_210 | _GEN_46; 
  assign _T_213 = _T_212[19:8]; 
  assign _GEN_47 = {{8'd0}, _T_213}; 
  assign _T_214 = _T_212 | _GEN_47; 
  assign _T_215 = _T_214[19:16]; 
  assign _GEN_48 = {{16'd0}, _T_215}; 
  assign _T_216 = _T_214 | _GEN_48; 
  assign _T_218 = _T_216[19:1]; 
  assign _T_219 = ~ rx_d; 
  assign _GEN_49 = {{1'd0}, _T_218}; 
  assign _T_220 = _T_219 | _GEN_49; 
  assign _T_221 = ~ _T_220; 
  assign _T_222 = {_T_221, 1'h0}; 
  assign _T_223 = _T_222[20:16]; 
  assign _T_224 = _T_222[15:0]; 
  assign _T_225 = _T_223 != 5'h0; 
  assign _GEN_50 = {{11'd0}, _T_223}; 
  assign _T_226 = _GEN_50 | _T_224; 
  assign _T_227 = _T_226[15:8]; 
  assign _T_228 = _T_226[7:0]; 
  assign _T_229 = _T_227 != 8'h0; 
  assign _T_230 = _T_227 | _T_228; 
  assign _T_231 = _T_230[7:4]; 
  assign _T_232 = _T_230[3:0]; 
  assign _T_233 = _T_231 != 4'h0; 
  assign _T_234 = _T_231 | _T_232; 
  assign _T_235 = _T_234[3:2]; 
  assign _T_236 = _T_234[1:0]; 
  assign _T_237 = _T_235 != 2'h0; 
  assign _T_238 = _T_235 | _T_236; 
  assign _T_239 = _T_238[1]; 
  assign rxLeft_d = rx_d & _GEN_49; 
  assign _T_247 = rx_e[19:1]; 
  assign _GEN_52 = {{1'd0}, _T_247}; 
  assign _T_248 = rx_e | _GEN_52; 
  assign _T_249 = _T_248[19:2]; 
  assign _GEN_53 = {{2'd0}, _T_249}; 
  assign _T_250 = _T_248 | _GEN_53; 
  assign _T_251 = _T_250[19:4]; 
  assign _GEN_54 = {{4'd0}, _T_251}; 
  assign _T_252 = _T_250 | _GEN_54; 
  assign _T_253 = _T_252[19:8]; 
  assign _GEN_55 = {{8'd0}, _T_253}; 
  assign _T_254 = _T_252 | _GEN_55; 
  assign _T_255 = _T_254[19:16]; 
  assign _GEN_56 = {{16'd0}, _T_255}; 
  assign _T_256 = _T_254 | _GEN_56; 
  assign _T_258 = _T_256[19:1]; 
  assign _T_259 = ~ rx_e; 
  assign _GEN_57 = {{1'd0}, _T_258}; 
  assign _T_260 = _T_259 | _GEN_57; 
  assign _T_261 = ~ _T_260; 
  assign _T_262 = {_T_261, 1'h0}; 
  assign _T_263 = _T_262[20:16]; 
  assign _T_264 = _T_262[15:0]; 
  assign _T_265 = _T_263 != 5'h0; 
  assign _GEN_58 = {{11'd0}, _T_263}; 
  assign _T_266 = _GEN_58 | _T_264; 
  assign _T_267 = _T_266[15:8]; 
  assign _T_268 = _T_266[7:0]; 
  assign _T_269 = _T_267 != 8'h0; 
  assign _T_270 = _T_267 | _T_268; 
  assign _T_271 = _T_270[7:4]; 
  assign _T_272 = _T_270[3:0]; 
  assign _T_273 = _T_271 != 4'h0; 
  assign _T_274 = _T_271 | _T_272; 
  assign _T_275 = _T_274[3:2]; 
  assign _T_276 = _T_274[1:0]; 
  assign _T_277 = _T_275 != 2'h0; 
  assign _T_278 = _T_275 | _T_276; 
  assign _T_279 = _T_278[1]; 
  assign rxLeft_e = rx_e & _GEN_57; 
  assign _T_288 = {_T_105,_T_109,_T_113,_T_117,_T_119,4'h0,3'h5}; 
  assign _T_289 = {_T_185,_T_189,_T_193,_T_197,_T_199,_T_145,_T_149,_T_153,_T_157,_T_159}; 
  assign _T_290 = {_T_265,_T_269,_T_273,_T_277,_T_279,_T_225,_T_229,_T_233,_T_237,_T_239}; 
  assign _T_291 = {_T_290,_T_289}; 
  assign _T_292 = rxQ_io_enq_ready & rxQ_io_enq_valid; 
  assign _T_293_a = _T_292 ? rxLeft_a : rx_a; 
  assign _T_293_b = _T_292 ? rxLeft_b : rx_b; 
  assign _T_293_c = _T_292 ? rxLeft_c : rx_c; 
  assign _T_293_d = _T_292 ? rxLeft_d : rx_d; 
  assign _T_293_e = _T_292 ? rxLeft_e : rx_e; 
  assign _T_294 = AsyncQueueSink_io_deq_ready & AsyncQueueSink_io_deq_valid; 
  assign _T_296_a = _T_294 ? AsyncQueueSink_io_deq_bits_a : 20'h0; 
  assign _T_296_b = _T_294 ? AsyncQueueSink_io_deq_bits_b : 20'h0; 
  assign _T_296_c = _T_294 ? AsyncQueueSink_io_deq_bits_c : 20'h0; 
  assign _T_296_d = _T_294 ? AsyncQueueSink_io_deq_bits_d : 20'h0; 
  assign _T_296_e = _T_294 ? AsyncQueueSink_io_deq_bits_e : 20'h0; 
  assign _T_298 = _T_293_a + _T_296_a; 
  assign _T_299 = _T_298[20:20]; 
  assign _T_302 = _T_299 ? 21'hfffff : _T_298; 
  assign _T_303 = _T_293_b + _T_296_b; 
  assign _T_304 = _T_303[20:20]; 
  assign _T_307 = _T_304 ? 21'hfffff : _T_303; 
  assign _T_308 = _T_293_c + _T_296_c; 
  assign _T_309 = _T_308[20:20]; 
  assign _T_312 = _T_309 ? 21'hfffff : _T_308; 
  assign _T_313 = _T_293_d + _T_296_d; 
  assign _T_314 = _T_313[20:20]; 
  assign _T_317 = _T_314 ? 21'hfffff : _T_313; 
  assign _T_318 = _T_293_e + _T_296_e; 
  assign _T_319 = _T_318[20:20]; 
  assign _T_322 = _T_319 ? 21'hfffff : _T_318; 
  assign _T_336 = ShiftQueue_5_io_deq_valid | ShiftQueue_6_io_deq_valid; 
  assign _T_337 = _T_336 | ShiftQueue_7_io_deq_valid; 
  assign _T_338 = _T_337 | ShiftQueue_8_io_deq_valid; 
  assign _T_339 = _T_338 | ShiftQueue_9_io_deq_valid; 
  assign _T_340 = _T_339 == 1'h0; 
  assign forceXmit = xmit == 5'h0; 
  assign allowReturn = _T_340 | forceXmit; 
  assign f_valid = rxQ_io_deq_valid & allowReturn; 
  assign requests = {f_valid,ShiftQueue_9_io_deq_valid,ShiftQueue_8_io_deq_valid,ShiftQueue_7_io_deq_valid,ShiftQueue_6_io_deq_valid,ShiftQueue_5_io_deq_valid}; 
  assign f_bits_last = rxQ_io_deq_bits_last; 
  assign lasts = {f_bits_last,ShiftQueue_9_io_deq_bits_last,ShiftQueue_8_io_deq_bits_last,ShiftQueue_7_io_deq_bits_last,ShiftQueue_6_io_deq_bits_last,ShiftQueue_5_io_deq_bits_last}; 
  assign _T_331 = forceXmit == 1'h0; 
  assign _T_333 = xmit - 5'h1; 
  assign _T_350 = ~ _T_349; 
  assign _T_351 = requests & _T_350; 
  assign _T_352 = {_T_351,f_valid,ShiftQueue_9_io_deq_valid,ShiftQueue_8_io_deq_valid,ShiftQueue_7_io_deq_valid,ShiftQueue_6_io_deq_valid,ShiftQueue_5_io_deq_valid}; 
  assign _T_353 = _T_352[11:1]; 
  assign _GEN_60 = {{1'd0}, _T_353}; 
  assign _T_354 = _T_352 | _GEN_60; 
  assign _T_355 = _T_354[11:2]; 
  assign _GEN_61 = {{2'd0}, _T_355}; 
  assign _T_356 = _T_354 | _GEN_61; 
  assign _T_357 = _T_356[11:4]; 
  assign _GEN_62 = {{4'd0}, _T_357}; 
  assign _T_358 = _T_356 | _GEN_62; 
  assign _T_360 = _T_358[11:1]; 
  assign _T_361 = {_T_349, 6'h0}; 
  assign _GEN_63 = {{1'd0}, _T_360}; 
  assign _T_362 = _GEN_63 | _T_361; 
  assign _T_363 = _T_362[11:6]; 
  assign _T_364 = _T_362[5:0]; 
  assign _T_365 = _T_363 & _T_364; 
  assign readys = ~ _T_365; 
  assign allowed = first ? readys : state; 
  assign f_ready = allowed[5]; 
  assign _T_334 = f_ready & f_valid; 
  assign _T_344 = requests == requests; 
  assign _T_346 = _T_344 | reset; 
  assign _T_347 = _T_346 == 1'h0; 
  assign _T_367 = requests != 6'h0; 
  assign _T_368 = first & _T_367; 
  assign _T_369 = readys & requests; 
  assign _T_370 = {_T_369, 1'h0}; 
  assign _T_371 = _T_370[5:0]; 
  assign _T_372 = _T_369 | _T_371; 
  assign _T_373 = {_T_372, 2'h0}; 
  assign _T_374 = _T_373[5:0]; 
  assign _T_375 = _T_372 | _T_374; 
  assign _T_376 = {_T_375, 4'h0}; 
  assign _T_377 = _T_376[5:0]; 
  assign _T_378 = _T_375 | _T_377; 
  assign grant = first ? _T_369 : state; 
  assign _T_386 = state & requests; 
  assign _T_387 = _T_386 != 6'h0; 
  assign send = first ? rxQ_io_deq_valid : _T_387; 
  assign _T_388 = grant & requests; 
  assign _T_389 = _T_388 != 6'h0; 
  assign _T_390 = send == _T_389; 
  assign _T_392 = _T_390 | reset; 
  assign _T_393 = _T_392 == 1'h0; 
  assign _T_394 = grant & lasts; 
  assign _T_395 = _T_394 != 6'h0; 
  assign _T_402 = _T_399[0]; 
  assign _T_403 = _T_399[1]; 
  assign _T_404 = _T_399[2]; 
  assign _T_405 = _T_399[3]; 
  assign _T_406 = _T_399[4]; 
  assign _T_407 = _T_399[5]; 
  assign _T_408 = _T_402 ? _T_401_0 : 32'h0; 
  assign _T_409 = _T_403 ? _T_401_1 : 32'h0; 
  assign _T_410 = _T_404 ? _T_401_2 : 32'h0; 
  assign _T_411 = _T_405 ? _T_401_3 : 32'h0; 
  assign _T_412 = _T_406 ? _T_401_4 : 32'h0; 
  assign _T_413 = _T_407 ? _T_401_5 : 32'h0; 
  assign _T_414 = _T_408 | _T_409; 
  assign _T_415 = _T_414 | _T_410; 
  assign _T_416 = _T_415 | _T_411; 
  assign _T_417 = _T_416 | _T_412; 
  assign _T_297_a = _T_302[19:0]; 
  assign _T_297_b = _T_307[19:0]; 
  assign _T_297_c = _T_312[19:0]; 
  assign _T_297_d = _T_317[19:0]; 
  assign _T_297_e = _T_322[19:0]; 
  assign io_c2b_clk = clock; 
  assign io_c2b_rst = AsyncResetReg_q; 
  assign io_c2b_send = _T_398; 
  assign io_c2b_data = _T_420; 
  assign io_sa_ready = ShiftQueue_io_enq_ready; 
  assign io_sb_ready = ShiftQueue_1_io_enq_ready; 
  assign io_sc_ready = ShiftQueue_2_io_enq_ready; 
  assign io_sd_ready = ShiftQueue_3_io_enq_ready; 
  assign io_rxc_ridx = AsyncQueueSink_io_async_ridx; 
  assign io_rxc_safe_ridx_valid = AsyncQueueSink_io_async_safe_ridx_valid; 
  assign io_rxc_safe_sink_reset_n = AsyncQueueSink_io_async_safe_sink_reset_n; 
  assign io_txc_ridx = AsyncQueueSink_1_io_async_ridx; 
  assign io_txc_safe_ridx_valid = AsyncQueueSink_1_io_async_safe_ridx_valid; 
  assign io_txc_safe_sink_reset_n = AsyncQueueSink_1_io_async_safe_sink_reset_n; 
  assign AsyncQueueSink_clock = clock; 
  assign AsyncQueueSink_reset = reset; 
  assign AsyncQueueSink_io_deq_ready = 1'h1; 
  assign AsyncQueueSink_io_async_mem_0_a = io_rxc_mem_0_a; 
  assign AsyncQueueSink_io_async_mem_0_b = io_rxc_mem_0_b; 
  assign AsyncQueueSink_io_async_mem_0_c = io_rxc_mem_0_c; 
  assign AsyncQueueSink_io_async_mem_0_d = io_rxc_mem_0_d; 
  assign AsyncQueueSink_io_async_mem_0_e = io_rxc_mem_0_e; 
  assign AsyncQueueSink_io_async_widx = io_rxc_widx; 
  assign AsyncQueueSink_io_async_safe_widx_valid = io_rxc_safe_widx_valid; 
  assign AsyncQueueSink_io_async_safe_source_reset_n = io_rxc_safe_source_reset_n; 
  assign AsyncQueueSink_1_clock = clock; 
  assign AsyncQueueSink_1_reset = reset; 
  assign AsyncQueueSink_1_io_deq_ready = 1'h1; 
  assign AsyncQueueSink_1_io_async_mem_0_a = io_txc_mem_0_a; 
  assign AsyncQueueSink_1_io_async_mem_0_b = io_txc_mem_0_b; 
  assign AsyncQueueSink_1_io_async_mem_0_c = io_txc_mem_0_c; 
  assign AsyncQueueSink_1_io_async_mem_0_d = io_txc_mem_0_d; 
  assign AsyncQueueSink_1_io_async_mem_0_e = io_txc_mem_0_e; 
  assign AsyncQueueSink_1_io_async_widx = io_txc_widx; 
  assign AsyncQueueSink_1_io_async_safe_widx_valid = io_txc_safe_widx_valid; 
  assign AsyncQueueSink_1_io_async_safe_source_reset_n = io_txc_safe_source_reset_n; 
  assign ShiftQueue_clock = clock; 
  assign ShiftQueue_reset = reset; 
  assign ShiftQueue_io_enq_valid = io_sa_valid; 
  assign ShiftQueue_io_enq_bits_data = io_sa_bits_data; 
  assign ShiftQueue_io_enq_bits_last = io_sa_bits_last; 
  assign ShiftQueue_io_enq_bits_beats = io_sa_bits_beats; 
  assign ShiftQueue_io_deq_ready = ShiftQueue_5_io_enq_ready & _T_9; 
  assign ShiftQueue_1_clock = clock; 
  assign ShiftQueue_1_reset = reset; 
  assign ShiftQueue_1_io_enq_valid = 1'h0; 
  assign ShiftQueue_1_io_enq_bits_data = io_sb_bits_data; 
  assign ShiftQueue_1_io_enq_bits_last = io_sb_bits_last; 
  assign ShiftQueue_1_io_enq_bits_beats = 13'h3; 
  assign ShiftQueue_1_io_deq_ready = ShiftQueue_6_io_enq_ready & _T_26; 
  assign ShiftQueue_2_clock = clock; 
  assign ShiftQueue_2_reset = reset; 
  assign ShiftQueue_2_io_enq_valid = 1'h0; 
  assign ShiftQueue_2_io_enq_bits_data = io_sc_bits_data; 
  assign ShiftQueue_2_io_enq_bits_last = io_sc_bits_last; 
  assign ShiftQueue_2_io_enq_bits_beats = 13'h3; 
  assign ShiftQueue_2_io_deq_ready = ShiftQueue_7_io_enq_ready & _T_43; 
  assign ShiftQueue_3_clock = clock; 
  assign ShiftQueue_3_reset = reset; 
  assign ShiftQueue_3_io_enq_valid = io_sd_valid; 
  assign ShiftQueue_3_io_enq_bits_data = io_sd_bits_data; 
  assign ShiftQueue_3_io_enq_bits_last = io_sd_bits_last; 
  assign ShiftQueue_3_io_enq_bits_beats = io_sd_bits_beats; 
  assign ShiftQueue_3_io_deq_ready = ShiftQueue_8_io_enq_ready & _T_60; 
  assign ShiftQueue_4_clock = clock; 
  assign ShiftQueue_4_reset = reset; 
  assign ShiftQueue_4_io_enq_valid = 1'h0; 
  assign ShiftQueue_4_io_enq_bits_data = io_se_bits_data; 
  assign ShiftQueue_4_io_enq_bits_last = 1'h1; 
  assign ShiftQueue_4_io_enq_bits_beats = 13'h1; 
  assign ShiftQueue_4_io_deq_ready = ShiftQueue_9_io_enq_ready & _T_77; 
  assign ShiftQueue_5_clock = clock; 
  assign ShiftQueue_5_reset = reset; 
  assign ShiftQueue_5_io_enq_valid = ShiftQueue_io_deq_valid & _T_9; 
  assign ShiftQueue_5_io_enq_bits_data = ShiftQueue_io_deq_bits_data; 
  assign ShiftQueue_5_io_enq_bits_last = ShiftQueue_io_deq_bits_last; 
  assign ShiftQueue_5_io_enq_bits_beats = ShiftQueue_io_deq_bits_beats; 
  assign ShiftQueue_5_io_deq_ready = allowed[0]; 
  assign ShiftQueue_6_clock = clock; 
  assign ShiftQueue_6_reset = reset; 
  assign ShiftQueue_6_io_enq_valid = ShiftQueue_1_io_deq_valid & _T_26; 
  assign ShiftQueue_6_io_enq_bits_data = ShiftQueue_1_io_deq_bits_data; 
  assign ShiftQueue_6_io_enq_bits_last = ShiftQueue_1_io_deq_bits_last; 
  assign ShiftQueue_6_io_enq_bits_beats = ShiftQueue_1_io_deq_bits_beats; 
  assign ShiftQueue_6_io_deq_ready = allowed[1]; 
  assign ShiftQueue_7_clock = clock; 
  assign ShiftQueue_7_reset = reset; 
  assign ShiftQueue_7_io_enq_valid = ShiftQueue_2_io_deq_valid & _T_43; 
  assign ShiftQueue_7_io_enq_bits_data = ShiftQueue_2_io_deq_bits_data; 
  assign ShiftQueue_7_io_enq_bits_last = ShiftQueue_2_io_deq_bits_last; 
  assign ShiftQueue_7_io_enq_bits_beats = ShiftQueue_2_io_deq_bits_beats; 
  assign ShiftQueue_7_io_deq_ready = allowed[2]; 
  assign ShiftQueue_8_clock = clock; 
  assign ShiftQueue_8_reset = reset; 
  assign ShiftQueue_8_io_enq_valid = ShiftQueue_3_io_deq_valid & _T_60; 
  assign ShiftQueue_8_io_enq_bits_data = ShiftQueue_3_io_deq_bits_data; 
  assign ShiftQueue_8_io_enq_bits_last = ShiftQueue_3_io_deq_bits_last; 
  assign ShiftQueue_8_io_enq_bits_beats = ShiftQueue_3_io_deq_bits_beats; 
  assign ShiftQueue_8_io_deq_ready = allowed[3]; 
  assign ShiftQueue_9_clock = clock; 
  assign ShiftQueue_9_reset = reset; 
  assign ShiftQueue_9_io_enq_valid = ShiftQueue_4_io_deq_valid & _T_77; 
  assign ShiftQueue_9_io_enq_bits_data = ShiftQueue_4_io_deq_bits_data; 
  assign ShiftQueue_9_io_enq_bits_last = ShiftQueue_4_io_deq_bits_last; 
  assign ShiftQueue_9_io_enq_bits_beats = ShiftQueue_4_io_deq_bits_beats; 
  assign ShiftQueue_9_io_deq_ready = allowed[4]; 
  assign rxQ_clock = clock; 
  assign rxQ_reset = reset; 
  assign rxQ_io_enq_valid = 1'h1; 
  assign rxQ_io_enq_bits_data = {_T_291,_T_288}; 
  assign rxQ_io_enq_bits_last = 1'h1; 
  assign rxQ_io_enq_bits_beats = 13'h1; 
  assign rxQ_io_deq_ready = f_ready & allowReturn; 
  assign AsyncResetReg_d = 1'h0; 
  assign AsyncResetReg_en = 1'h1; 
  assign AsyncResetReg_clk = clock; 
  assign AsyncResetReg_rst = reset; 
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rx_a = _RAND_0[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  rx_b = _RAND_1[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  rx_c = _RAND_2[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  rx_d = _RAND_3[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  rx_e = _RAND_4[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  tx_a = _RAND_5[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  tx_b = _RAND_6[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  tx_c = _RAND_7[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  tx_d = _RAND_8[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  tx_e = _RAND_9[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_3 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_20 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_37 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_54 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_71 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  xmit = _RAND_15[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  first = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_349 = _RAND_17[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  state = _RAND_18[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_397 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_398 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_399 = _RAND_21[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_401_0 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_401_1 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_401_2 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_401_3 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_401_4 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_401_5 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_420 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      rx_a <= 20'h0;
    end else begin
      rx_a <= _T_297_a;
    end
    if (reset) begin
      rx_b <= 20'h0;
    end else begin
      rx_b <= _T_297_b;
    end
    if (reset) begin
      rx_c <= 20'h0;
    end else begin
      rx_c <= _T_297_c;
    end
    if (reset) begin
      rx_d <= 20'h0;
    end else begin
      rx_d <= _T_297_d;
    end
    if (reset) begin
      rx_e <= 20'h0;
    end else begin
      rx_e <= _T_297_e;
    end
    if (reset) begin
      tx_a <= 20'h0;
    end else begin
      tx_a <= _T_16[19:0];
    end
    if (reset) begin
      tx_b <= 20'h0;
    end else begin
      tx_b <= _T_33[19:0];
    end
    if (reset) begin
      tx_c <= 20'h0;
    end else begin
      tx_c <= _T_50[19:0];
    end
    if (reset) begin
      tx_d <= 20'h0;
    end else begin
      tx_d <= _T_67[19:0];
    end
    if (reset) begin
      tx_e <= 20'h0;
    end else begin
      tx_e <= _T_84[19:0];
    end
    if (reset) begin
      _T_3 <= 1'h1;
    end else begin
      if (_T_2) begin
        _T_3 <= ShiftQueue_io_deq_bits_last;
      end
    end
    if (reset) begin
      _T_20 <= 1'h1;
    end else begin
      if (_T_19) begin
        _T_20 <= ShiftQueue_1_io_deq_bits_last;
      end
    end
    if (reset) begin
      _T_37 <= 1'h1;
    end else begin
      if (_T_36) begin
        _T_37 <= ShiftQueue_2_io_deq_bits_last;
      end
    end
    if (reset) begin
      _T_54 <= 1'h1;
    end else begin
      if (_T_53) begin
        _T_54 <= ShiftQueue_3_io_deq_bits_last;
      end
    end
    if (reset) begin
      _T_71 <= 1'h1;
    end else begin
      if (_T_70) begin
        _T_71 <= ShiftQueue_4_io_deq_bits_last;
      end
    end
    if (reset) begin
      xmit <= 5'h0;
    end else begin
      if (_T_334) begin
        xmit <= 5'h1f;
      end else begin
        if (_T_331) begin
          xmit <= _T_333;
        end
      end
    end
    if (reset) begin
      first <= 1'h1;
    end else begin
      if (send) begin
        first <= _T_395;
      end
    end
    if (reset) begin
      _T_349 <= 6'h3f;
    end else begin
      if (_T_368) begin
        _T_349 <= _T_378;
      end
    end
    if (first) begin
      state <= _T_369;
    end
    if (reset) begin
      _T_397 <= 1'h0;
    end else begin
      if (first) begin
        _T_397 <= rxQ_io_deq_valid;
      end else begin
        _T_397 <= _T_387;
      end
    end
    if (reset) begin
      _T_398 <= 1'h0;
    end else begin
      _T_398 <= _T_397;
    end
    if (first) begin
      _T_399 <= _T_369;
    end else begin
      _T_399 <= state;
    end
    _T_401_0 <= ShiftQueue_5_io_deq_bits_data;
    _T_401_1 <= ShiftQueue_6_io_deq_bits_data;
    _T_401_2 <= ShiftQueue_7_io_deq_bits_data;
    _T_401_3 <= ShiftQueue_8_io_deq_bits_data;
    _T_401_4 <= ShiftQueue_9_io_deq_bits_data;
    _T_401_5 <= rxQ_io_deq_bits_data;
    _T_420 <= _T_417 | _T_413;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_347) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_347) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_393) begin
          $fwrite(32'h80000002,"Assertion failed\n    at dual_TX.scala:100 assert (send === ((grant & requests) =/= UInt(0)))\n"); 
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_393) begin
          $fatal; 
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
